
module Midori64Enc ( clk, rst, Plaintext, Key, Ciphertext, done );
  input [63:0] Plaintext;
  input [127:0] Key;
  output [63:0] Ciphertext;
  input clk, rst;
  output done;
  wire   FSM[4] , AddKeyConstXOR_XORInst_0_0_N1 ,
         AddKeyConstXOR_XORInst_0_1_N0 , AddKeyConstXOR_XORInst_0_2_N0 ,
         AddKeyConstXOR_XORInst_0_3_N0 , AddKeyConstXOR_XORInst_1_0_N1 ,
         AddKeyConstXOR_XORInst_1_1_N0 , AddKeyConstXOR_XORInst_1_2_N0 ,
         AddKeyConstXOR_XORInst_1_3_N0 , AddKeyConstXOR_XORInst_2_0_N1 ,
         AddKeyConstXOR_XORInst_2_1_N0 , AddKeyConstXOR_XORInst_2_2_N0 ,
         AddKeyConstXOR_XORInst_2_3_N0 , AddKeyConstXOR_XORInst_3_0_N1 ,
         AddKeyConstXOR_XORInst_3_1_N0 , AddKeyConstXOR_XORInst_3_2_N0 ,
         AddKeyConstXOR_XORInst_3_3_N0 , AddKeyConstXOR_XORInst_4_0_N1 ,
         AddKeyConstXOR_XORInst_4_1_N0 , AddKeyConstXOR_XORInst_4_2_N0 ,
         AddKeyConstXOR_XORInst_4_3_N0 , AddKeyConstXOR_XORInst_5_0_N1 ,
         AddKeyConstXOR_XORInst_5_1_N0 , AddKeyConstXOR_XORInst_5_2_N0 ,
         AddKeyConstXOR_XORInst_5_3_N0 , AddKeyConstXOR_XORInst_6_0_N1 ,
         AddKeyConstXOR_XORInst_6_1_N0 , AddKeyConstXOR_XORInst_6_2_N0 ,
         AddKeyConstXOR_XORInst_6_3_N0 , AddKeyConstXOR_XORInst_7_0_N1 ,
         AddKeyConstXOR_XORInst_7_1_N0 , AddKeyConstXOR_XORInst_7_2_N0 ,
         AddKeyConstXOR_XORInst_7_3_N0 , AddKeyConstXOR_XORInst_8_0_N1 ,
         AddKeyConstXOR_XORInst_8_1_N0 , AddKeyConstXOR_XORInst_8_2_N0 ,
         AddKeyConstXOR_XORInst_8_3_N0 , AddKeyConstXOR_XORInst_9_0_N1 ,
         AddKeyConstXOR_XORInst_9_1_N0 , AddKeyConstXOR_XORInst_9_2_N0 ,
         AddKeyConstXOR_XORInst_9_3_N0 , AddKeyConstXOR_XORInst_10_0_N1 ,
         AddKeyConstXOR_XORInst_10_1_N0 , AddKeyConstXOR_XORInst_10_2_N0 ,
         AddKeyConstXOR_XORInst_10_3_N0 , AddKeyConstXOR_XORInst_11_0_N1 ,
         AddKeyConstXOR_XORInst_11_1_N0 , AddKeyConstXOR_XORInst_11_2_N0 ,
         AddKeyConstXOR_XORInst_11_3_N0 , AddKeyConstXOR_XORInst_12_0_N1 ,
         AddKeyConstXOR_XORInst_12_1_N0 , AddKeyConstXOR_XORInst_12_2_N0 ,
         AddKeyConstXOR_XORInst_12_3_N0 , AddKeyConstXOR_XORInst_13_0_N1 ,
         AddKeyConstXOR_XORInst_13_1_N0 , AddKeyConstXOR_XORInst_13_2_N0 ,
         AddKeyConstXOR_XORInst_13_3_N0 , AddKeyConstXOR_XORInst_14_0_N1 ,
         AddKeyConstXOR_XORInst_14_1_N0 , AddKeyConstXOR_XORInst_14_2_N0 ,
         AddKeyConstXOR_XORInst_14_3_N0 , AddKeyConstXOR_XORInst_15_0_N1 ,
         AddKeyConstXOR_XORInst_15_1_N0 , AddKeyConstXOR_XORInst_15_2_N0 ,
         AddKeyConstXOR_XORInst_15_3_N0 , n1245, n1246, n1247, n1248, n1249,
         n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259,
         n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269,
         n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279,
         n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289,
         n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299,
         n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309,
         n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319,
         n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409,
         n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419,
         n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429,
         n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439,
         n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449,
         n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459,
         n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469,
         n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479,
         n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489,
         n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499,
         n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509,
         n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519,
         n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529,
         n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539,
         n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549,
         n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559,
         n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569,
         n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579,
         n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728, n1729,
         n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738, n1739,
         n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748, n1749,
         n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758, n1759,
         n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768, n1769,
         n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778, n1779,
         n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788, n1789,
         n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798, n1799,
         n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808, n1809,
         n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818, n1819,
         n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828, n1829,
         n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838, n1839,
         n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848, n1849,
         n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858, n1859,
         n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869,
         n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1879,
         n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888, n1889,
         n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898, n1899,
         n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908, n1909,
         n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918, n1919,
         n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928, n1929,
         n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938, n1939,
         n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948, n1949,
         n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958, n1959,
         n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968, n1969,
         n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978, n1979,
         n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988, n1989,
         n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998, n1999,
         n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008, n2009,
         n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018, n2019,
         n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028, n2029,
         n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038, n2039,
         n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048, n2049,
         n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058, n2059,
         n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068, n2069,
         n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078, n2079,
         n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088, n2089,
         n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098, n2099,
         n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108, n2109,
         n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118, n2119,
         n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128, n2129,
         n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138, n2139,
         n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148, n2149,
         n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158, n2159,
         n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168, n2169,
         n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178, n2179,
         n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188, n2189,
         n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198, n2199,
         n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208, n2209,
         n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218, n2219,
         n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228, n2229,
         n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238, n2239,
         n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248, n2249,
         n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258, n2259,
         n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268, n2269,
         n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278, n2279,
         n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288, n2289,
         n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298, n2299,
         n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308, n2309,
         n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318, n2319,
         n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328, n2329,
         n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338, n2339,
         n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348, n2349,
         n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358, n2359,
         n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368, n2369,
         n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378, n2379,
         n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388, n2389,
         n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398, n2399,
         n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408, n2409,
         n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418, n2419,
         n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428, n2429,
         n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438, n2439,
         n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448, n2449,
         n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458, n2459,
         n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468, n2469,
         n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478, n2479,
         n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488, n2489,
         n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498, n2499,
         n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508, n2509,
         n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518, n2519,
         n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528, n2529,
         n2530, n2531, n2532, n2533, n2534, n2535, n2536;
  wire   [63:0] StateRegInput;
  wire   [63:0] StateRegOutput;
  wire   [3:0] Round;
  wire   [4:0] FSMSelected;
  assign Ciphertext[0] = AddKeyConstXOR_XORInst_0_0_N1 ;
  assign Ciphertext[1] = AddKeyConstXOR_XORInst_0_1_N0 ;
  assign Ciphertext[2] = AddKeyConstXOR_XORInst_0_2_N0 ;
  assign Ciphertext[3] = AddKeyConstXOR_XORInst_0_3_N0 ;
  assign Ciphertext[4] = AddKeyConstXOR_XORInst_1_0_N1 ;
  assign Ciphertext[5] = AddKeyConstXOR_XORInst_1_1_N0 ;
  assign Ciphertext[6] = AddKeyConstXOR_XORInst_1_2_N0 ;
  assign Ciphertext[7] = AddKeyConstXOR_XORInst_1_3_N0 ;
  assign Ciphertext[8] = AddKeyConstXOR_XORInst_2_0_N1 ;
  assign Ciphertext[9] = AddKeyConstXOR_XORInst_2_1_N0 ;
  assign Ciphertext[10] = AddKeyConstXOR_XORInst_2_2_N0 ;
  assign Ciphertext[11] = AddKeyConstXOR_XORInst_2_3_N0 ;
  assign Ciphertext[12] = AddKeyConstXOR_XORInst_3_0_N1 ;
  assign Ciphertext[13] = AddKeyConstXOR_XORInst_3_1_N0 ;
  assign Ciphertext[14] = AddKeyConstXOR_XORInst_3_2_N0 ;
  assign Ciphertext[15] = AddKeyConstXOR_XORInst_3_3_N0 ;
  assign Ciphertext[16] = AddKeyConstXOR_XORInst_4_0_N1 ;
  assign Ciphertext[17] = AddKeyConstXOR_XORInst_4_1_N0 ;
  assign Ciphertext[18] = AddKeyConstXOR_XORInst_4_2_N0 ;
  assign Ciphertext[19] = AddKeyConstXOR_XORInst_4_3_N0 ;
  assign Ciphertext[20] = AddKeyConstXOR_XORInst_5_0_N1 ;
  assign Ciphertext[21] = AddKeyConstXOR_XORInst_5_1_N0 ;
  assign Ciphertext[22] = AddKeyConstXOR_XORInst_5_2_N0 ;
  assign Ciphertext[23] = AddKeyConstXOR_XORInst_5_3_N0 ;
  assign Ciphertext[24] = AddKeyConstXOR_XORInst_6_0_N1 ;
  assign Ciphertext[25] = AddKeyConstXOR_XORInst_6_1_N0 ;
  assign Ciphertext[26] = AddKeyConstXOR_XORInst_6_2_N0 ;
  assign Ciphertext[27] = AddKeyConstXOR_XORInst_6_3_N0 ;
  assign Ciphertext[28] = AddKeyConstXOR_XORInst_7_0_N1 ;
  assign Ciphertext[29] = AddKeyConstXOR_XORInst_7_1_N0 ;
  assign Ciphertext[30] = AddKeyConstXOR_XORInst_7_2_N0 ;
  assign Ciphertext[31] = AddKeyConstXOR_XORInst_7_3_N0 ;
  assign Ciphertext[32] = AddKeyConstXOR_XORInst_8_0_N1 ;
  assign Ciphertext[33] = AddKeyConstXOR_XORInst_8_1_N0 ;
  assign Ciphertext[34] = AddKeyConstXOR_XORInst_8_2_N0 ;
  assign Ciphertext[35] = AddKeyConstXOR_XORInst_8_3_N0 ;
  assign Ciphertext[36] = AddKeyConstXOR_XORInst_9_0_N1 ;
  assign Ciphertext[37] = AddKeyConstXOR_XORInst_9_1_N0 ;
  assign Ciphertext[38] = AddKeyConstXOR_XORInst_9_2_N0 ;
  assign Ciphertext[39] = AddKeyConstXOR_XORInst_9_3_N0 ;
  assign Ciphertext[40] = AddKeyConstXOR_XORInst_10_0_N1 ;
  assign Ciphertext[41] = AddKeyConstXOR_XORInst_10_1_N0 ;
  assign Ciphertext[42] = AddKeyConstXOR_XORInst_10_2_N0 ;
  assign Ciphertext[43] = AddKeyConstXOR_XORInst_10_3_N0 ;
  assign Ciphertext[44] = AddKeyConstXOR_XORInst_11_0_N1 ;
  assign Ciphertext[45] = AddKeyConstXOR_XORInst_11_1_N0 ;
  assign Ciphertext[46] = AddKeyConstXOR_XORInst_11_2_N0 ;
  assign Ciphertext[47] = AddKeyConstXOR_XORInst_11_3_N0 ;
  assign Ciphertext[48] = AddKeyConstXOR_XORInst_12_0_N1 ;
  assign Ciphertext[49] = AddKeyConstXOR_XORInst_12_1_N0 ;
  assign Ciphertext[50] = AddKeyConstXOR_XORInst_12_2_N0 ;
  assign Ciphertext[51] = AddKeyConstXOR_XORInst_12_3_N0 ;
  assign Ciphertext[52] = AddKeyConstXOR_XORInst_13_0_N1 ;
  assign Ciphertext[53] = AddKeyConstXOR_XORInst_13_1_N0 ;
  assign Ciphertext[54] = AddKeyConstXOR_XORInst_13_2_N0 ;
  assign Ciphertext[55] = AddKeyConstXOR_XORInst_13_3_N0 ;
  assign Ciphertext[56] = AddKeyConstXOR_XORInst_14_0_N1 ;
  assign Ciphertext[57] = AddKeyConstXOR_XORInst_14_1_N0 ;
  assign Ciphertext[58] = AddKeyConstXOR_XORInst_14_2_N0 ;
  assign Ciphertext[59] = AddKeyConstXOR_XORInst_14_3_N0 ;
  assign Ciphertext[60] = AddKeyConstXOR_XORInst_15_0_N1 ;
  assign Ciphertext[61] = AddKeyConstXOR_XORInst_15_1_N0 ;
  assign Ciphertext[62] = AddKeyConstXOR_XORInst_15_2_N0 ;
  assign Ciphertext[63] = AddKeyConstXOR_XORInst_15_3_N0 ;

  DFF FSMReg_s_current_state_reg[4]  ( .D(FSMSelected[4]), .CP(clk), .Q(
        FSM[4] ) );
  DFF FSMReg_s_current_state_reg[2]  ( .D(FSMSelected[2]), .CP(clk), .Q(
        Round[2]) );
  DFF FSMReg_s_current_state_reg[1]  ( .D(FSMSelected[1]), .CP(clk), .Q(
        Round[1]) );
  DFF FSMReg_s_current_state_reg[0]  ( .D(FSMSelected[0]), .CP(clk), .Q(
        Round[0]) );
  DFF FSMReg_s_current_state_reg[3]  ( .D(FSMSelected[3]), .CP(clk), .Q(
        Round[3]) );
  DFF StateReg_s_current_state_reg[13]  ( .D(StateRegInput[13]), .CP(clk), 
        .Q(StateRegOutput[13]) );
  DFF StateReg_s_current_state_reg[31]  ( .D(StateRegInput[31]), .CP(clk), 
        .Q(StateRegOutput[31]) );
  DFF StateReg_s_current_state_reg[29]  ( .D(StateRegInput[29]), .CP(clk), 
        .Q(StateRegOutput[29]) );
  DFF StateReg_s_current_state_reg[12]  ( .D(StateRegInput[12]), .CP(clk), 
        .Q(StateRegOutput[12]) );
  DFF StateReg_s_current_state_reg[14]  ( .D(StateRegInput[14]), .CP(clk), 
        .Q(StateRegOutput[14]) );
  DFF StateReg_s_current_state_reg[17]  ( .D(StateRegInput[17]), .CP(clk), 
        .Q(StateRegOutput[17]) );
  DFF StateReg_s_current_state_reg[19]  ( .D(StateRegInput[19]), .CP(clk), 
        .Q(StateRegOutput[19]) );
  DFF StateReg_s_current_state_reg[18]  ( .D(StateRegInput[18]), .CP(clk), 
        .Q(StateRegOutput[18]) );
  DFF StateReg_s_current_state_reg[33]  ( .D(StateRegInput[33]), .CP(clk), 
        .Q(StateRegOutput[33]) );
  DFF StateReg_s_current_state_reg[11]  ( .D(StateRegInput[11]), .CP(clk), 
        .Q(StateRegOutput[11]) );
  DFF StateReg_s_current_state_reg[1]  ( .D(StateRegInput[1]), .CP(clk), .Q(
        StateRegOutput[1]) );
  DFF StateReg_s_current_state_reg[63]  ( .D(StateRegInput[63]), .CP(clk), 
        .Q(StateRegOutput[63]) );
  DFF StateReg_s_current_state_reg[50]  ( .D(StateRegInput[50]), .CP(clk), 
        .Q(StateRegOutput[50]) );
  DFF StateReg_s_current_state_reg[21]  ( .D(StateRegInput[21]), .CP(clk), 
        .Q(StateRegOutput[21]) );
  DFF StateReg_s_current_state_reg[23]  ( .D(StateRegInput[23]), .CP(clk), 
        .Q(StateRegOutput[23]) );
  DFF StateReg_s_current_state_reg[22]  ( .D(StateRegInput[22]), .CP(clk), 
        .Q(StateRegOutput[22]) );
  DFF StateReg_s_current_state_reg[49]  ( .D(StateRegInput[49]), .CP(clk), 
        .Q(StateRegOutput[49]) );
  DFF StateReg_s_current_state_reg[51]  ( .D(StateRegInput[51]), .CP(clk), 
        .Q(StateRegOutput[51]) );
  DFF StateReg_s_current_state_reg[30]  ( .D(StateRegInput[30]), .CP(clk), 
        .Q(StateRegOutput[30]) );
  DFF StateReg_s_current_state_reg[15]  ( .D(StateRegInput[15]), .CP(clk), 
        .Q(StateRegOutput[15]) );
  DFF StateReg_s_current_state_reg[16]  ( .D(StateRegInput[16]), .CP(clk), 
        .Q(StateRegOutput[16]) );
  DFF StateReg_s_current_state_reg[32]  ( .D(StateRegInput[32]), .CP(clk), 
        .Q(StateRegOutput[32]) );
  DFF StateReg_s_current_state_reg[9]  ( .D(StateRegInput[9]), .CP(clk), .Q(
        StateRegOutput[9]) );
  DFF StateReg_s_current_state_reg[3]  ( .D(StateRegInput[3]), .CP(clk), .Q(
        StateRegOutput[3]) );
  DFF StateReg_s_current_state_reg[2]  ( .D(StateRegInput[2]), .CP(clk), .Q(
        StateRegOutput[2]) );
  DFF StateReg_s_current_state_reg[53]  ( .D(StateRegInput[53]), .CP(clk), 
        .Q(StateRegOutput[53]) );
  DFF StateReg_s_current_state_reg[55]  ( .D(StateRegInput[55]), .CP(clk), 
        .Q(StateRegOutput[55]) );
  DFF StateReg_s_current_state_reg[54]  ( .D(StateRegInput[54]), .CP(clk), 
        .Q(StateRegOutput[54]) );
  DFF StateReg_s_current_state_reg[10]  ( .D(StateRegInput[10]), .CP(clk), 
        .Q(StateRegOutput[10]) );
  DFF StateReg_s_current_state_reg[6]  ( .D(StateRegInput[6]), .CP(clk), .Q(
        StateRegOutput[6]) );
  DFF StateReg_s_current_state_reg[5]  ( .D(StateRegInput[5]), .CP(clk), .Q(
        StateRegOutput[5]) );
  DFF StateReg_s_current_state_reg[37]  ( .D(StateRegInput[37]), .CP(clk), 
        .Q(StateRegOutput[37]) );
  DFF StateReg_s_current_state_reg[27]  ( .D(StateRegInput[27]), .CP(clk), 
        .Q(StateRegOutput[27]) );
  DFF StateReg_s_current_state_reg[26]  ( .D(StateRegInput[26]), .CP(clk), 
        .Q(StateRegOutput[26]) );
  DFF StateReg_s_current_state_reg[25]  ( .D(StateRegInput[25]), .CP(clk), 
        .Q(StateRegOutput[25]) );
  DFF StateReg_s_current_state_reg[20]  ( .D(StateRegInput[20]), .CP(clk), 
        .Q(StateRegOutput[20]) );
  DFF StateReg_s_current_state_reg[60]  ( .D(StateRegInput[60]), .CP(clk), 
        .Q(StateRegOutput[60]) );
  DFF StateReg_s_current_state_reg[59]  ( .D(StateRegInput[59]), .CP(clk), 
        .Q(StateRegOutput[59]) );
  DFF StateReg_s_current_state_reg[42]  ( .D(StateRegInput[42]), .CP(clk), 
        .Q(StateRegOutput[42]) );
  DFF StateReg_s_current_state_reg[41]  ( .D(StateRegInput[41]), .CP(clk), 
        .Q(StateRegOutput[41]) );
  DFF StateReg_s_current_state_reg[43]  ( .D(StateRegInput[43]), .CP(clk), 
        .Q(StateRegOutput[43]) );
  DFF StateReg_s_current_state_reg[62]  ( .D(StateRegInput[62]), .CP(clk), 
        .Q(StateRegOutput[62]) );
  DFF StateReg_s_current_state_reg[61]  ( .D(StateRegInput[61]), .CP(clk), 
        .Q(StateRegOutput[61]) );
  DFF StateReg_s_current_state_reg[58]  ( .D(StateRegInput[58]), .CP(clk), 
        .Q(StateRegOutput[58]) );
  DFF StateReg_s_current_state_reg[57]  ( .D(StateRegInput[57]), .CP(clk), 
        .Q(StateRegOutput[57]) );
  DFF StateReg_s_current_state_reg[45]  ( .D(StateRegInput[45]), .CP(clk), 
        .Q(StateRegOutput[45]) );
  DFF StateReg_s_current_state_reg[35]  ( .D(StateRegInput[35]), .CP(clk), 
        .Q(StateRegOutput[35]) );
  DFF StateReg_s_current_state_reg[34]  ( .D(StateRegInput[34]), .CP(clk), 
        .Q(StateRegOutput[34]) );
  DFF StateReg_s_current_state_reg[8]  ( .D(StateRegInput[8]), .CP(clk), .Q(
        StateRegOutput[8]) );
  DFF StateReg_s_current_state_reg[4]  ( .D(StateRegInput[4]), .CP(clk), .Q(
        StateRegOutput[4]) );
  DFF StateReg_s_current_state_reg[7]  ( .D(StateRegInput[7]), .CP(clk), .Q(
        StateRegOutput[7]) );
  DFF StateReg_s_current_state_reg[0]  ( .D(StateRegInput[0]), .CP(clk), .Q(
        StateRegOutput[0]) );
  DFF StateReg_s_current_state_reg[56]  ( .D(StateRegInput[56]), .CP(clk), 
        .Q(StateRegOutput[56]) );
  DFF StateReg_s_current_state_reg[40]  ( .D(StateRegInput[40]), .CP(clk), 
        .Q(StateRegOutput[40]) );
  DFF StateReg_s_current_state_reg[39]  ( .D(StateRegInput[39]), .CP(clk), 
        .Q(StateRegOutput[39]) );
  DFF StateReg_s_current_state_reg[47]  ( .D(StateRegInput[47]), .CP(clk), 
        .Q(StateRegOutput[47]) );
  DFF StateReg_s_current_state_reg[46]  ( .D(StateRegInput[46]), .CP(clk), 
        .Q(StateRegOutput[46]) );
  DFF StateReg_s_current_state_reg[44]  ( .D(StateRegInput[44]), .CP(clk), 
        .Q(StateRegOutput[44]) );
  DFF StateReg_s_current_state_reg[38]  ( .D(StateRegInput[38]), .CP(clk), 
        .Q(StateRegOutput[38]) );
  DFF StateReg_s_current_state_reg[36]  ( .D(StateRegInput[36]), .CP(clk), 
        .Q(StateRegOutput[36]) );
  DFF StateReg_s_current_state_reg[24]  ( .D(StateRegInput[24]), .CP(clk), 
        .Q(StateRegOutput[24]) );
  DFF StateReg_s_current_state_reg[52]  ( .D(StateRegInput[52]), .CP(clk), 
        .Q(StateRegOutput[52]) );
  DFF StateReg_s_current_state_reg[48]  ( .D(StateRegInput[48]), .CP(clk), 
        .Q(StateRegOutput[48]) );
  DFF StateReg_s_current_state_reg[28]  ( .D(StateRegInput[28]), .CP(clk), 
        .Q(StateRegOutput[28]) );
  BIC2 U1380 ( .A(FSM[4] ), .B(Round[0]), .Z(done) );
  ORN2 U1381 ( .A(n1245), .B(n1246), .Z(StateRegInput[9]) );
  AND2 U1382 ( .A(n1247), .B(n1248), .Z(n1246) );
  ORN2 U1383 ( .A(n1249), .B(n1250), .Z(n1248) );
  XOR2 U1384 ( .A(n1251), .B(n1252), .Z(n1250) );
  NOT1 U1385 ( .A(n1253), .Z(n1252) );
  ORN2 U1386 ( .A(n1254), .B(n1255), .Z(n1247) );
  AND2 U1387 ( .A(Plaintext[9]), .B(rst), .Z(n1245) );
  ORN2 U1388 ( .A(n1256), .B(n1257), .Z(StateRegInput[8]) );
  AND2 U1389 ( .A(n1258), .B(n1259), .Z(n1257) );
  ORN2 U1390 ( .A(n1260), .B(n1261), .Z(n1259) );
  XOR2 U1391 ( .A(n1262), .B(n1263), .Z(n1260) );
  ORN2 U1392 ( .A(n1254), .B(n1264), .Z(n1258) );
  AND2 U1393 ( .A(Plaintext[8]), .B(rst), .Z(n1256) );
  ORN2 U1394 ( .A(n1265), .B(n1266), .Z(StateRegInput[7]) );
  AND2 U1395 ( .A(n1267), .B(n1268), .Z(n1266) );
  ORN2 U1396 ( .A(n1269), .B(n1261), .Z(n1268) );
  XOR2 U1397 ( .A(n1270), .B(n1271), .Z(n1269) );
  ORN2 U1398 ( .A(n1272), .B(n1273), .Z(n1267) );
  AND2 U1399 ( .A(Plaintext[7]), .B(rst), .Z(n1265) );
  ORN2 U1400 ( .A(n1274), .B(n1275), .Z(StateRegInput[6]) );
  AND2 U1401 ( .A(n1276), .B(n1277), .Z(n1275) );
  ORN2 U1402 ( .A(n1278), .B(n1261), .Z(n1277) );
  XOR2 U1403 ( .A(n1279), .B(n1280), .Z(n1278) );
  ORN2 U1404 ( .A(n1281), .B(n1273), .Z(n1276) );
  AND2 U1405 ( .A(Plaintext[6]), .B(rst), .Z(n1274) );
  ORN2 U1406 ( .A(n1282), .B(n1283), .Z(StateRegInput[63]) );
  AND2 U1407 ( .A(n1284), .B(n1285), .Z(n1283) );
  ORN2 U1408 ( .A(n1249), .B(n1286), .Z(n1285) );
  XOR2 U1409 ( .A(n1287), .B(n1288), .Z(n1286) );
  ORN2 U1410 ( .A(n1254), .B(n1289), .Z(n1284) );
  AND2 U1411 ( .A(Plaintext[63]), .B(rst), .Z(n1282) );
  ORN2 U1412 ( .A(n1290), .B(n1291), .Z(StateRegInput[62]) );
  AND2 U1413 ( .A(n1292), .B(n1293), .Z(n1291) );
  ORN2 U1414 ( .A(n1294), .B(n1261), .Z(n1293) );
  XOR2 U1415 ( .A(n1295), .B(n1296), .Z(n1294) );
  ORN2 U1416 ( .A(n1254), .B(n1297), .Z(n1292) );
  AND2 U1417 ( .A(Plaintext[62]), .B(rst), .Z(n1290) );
  ORN2 U1418 ( .A(n1298), .B(n1299), .Z(StateRegInput[61]) );
  AND2 U1419 ( .A(n1300), .B(n1301), .Z(n1299) );
  ORN2 U1420 ( .A(n1249), .B(n1302), .Z(n1301) );
  XOR2 U1421 ( .A(n1303), .B(n1304), .Z(n1302) );
  ORN2 U1422 ( .A(n1254), .B(n1305), .Z(n1300) );
  AND2 U1423 ( .A(Plaintext[61]), .B(rst), .Z(n1298) );
  ORN2 U1424 ( .A(n1306), .B(n1307), .Z(StateRegInput[60]) );
  AND2 U1425 ( .A(n1308), .B(n1309), .Z(n1307) );
  ORN2 U1426 ( .A(n1310), .B(n1261), .Z(n1309) );
  XOR2 U1427 ( .A(n1311), .B(n1312), .Z(n1310) );
  ORN2 U1428 ( .A(n1254), .B(n1313), .Z(n1308) );
  AND2 U1429 ( .A(Plaintext[60]), .B(rst), .Z(n1306) );
  ORN2 U1430 ( .A(n1314), .B(n1315), .Z(StateRegInput[5]) );
  AND2 U1431 ( .A(n1316), .B(n1317), .Z(n1315) );
  ORN2 U1432 ( .A(n1249), .B(n1318), .Z(n1317) );
  XOR2 U1433 ( .A(n1319), .B(n1320), .Z(n1318) );
  ORN2 U1434 ( .A(n1254), .B(n1321), .Z(n1316) );
  AND2 U1435 ( .A(Plaintext[5]), .B(rst), .Z(n1314) );
  ORN2 U1436 ( .A(n1322), .B(n1323), .Z(StateRegInput[59]) );
  AND2 U1437 ( .A(n1324), .B(n1325), .Z(n1323) );
  ORN2 U1438 ( .A(n1326), .B(n1261), .Z(n1325) );
  XOR2 U1439 ( .A(n1287), .B(n1289), .Z(n1326) );
  XOR2 U1440 ( .A(n1327), .B(n1328), .Z(n1287) );
  ORN2 U1441 ( .A(n1254), .B(n1329), .Z(n1324) );
  AND2 U1442 ( .A(Plaintext[59]), .B(rst), .Z(n1322) );
  ORN2 U1443 ( .A(n1330), .B(n1331), .Z(StateRegInput[58]) );
  AND2 U1444 ( .A(n1332), .B(n1333), .Z(n1331) );
  ORN2 U1445 ( .A(n1249), .B(n1334), .Z(n1333) );
  XOR2 U1446 ( .A(n1295), .B(n1297), .Z(n1334) );
  XOR2 U1447 ( .A(n1335), .B(n1336), .Z(n1295) );
  ORN2 U1448 ( .A(n1337), .B(n1273), .Z(n1332) );
  AND2 U1449 ( .A(Plaintext[58]), .B(rst), .Z(n1330) );
  ORN2 U1450 ( .A(n1338), .B(n1339), .Z(StateRegInput[57]) );
  AND2 U1451 ( .A(n1340), .B(n1341), .Z(n1339) );
  OR2 U1452 ( .A(n1342), .B(n1249), .Z(n1341) );
  XOR2 U1453 ( .A(n1303), .B(n1305), .Z(n1342) );
  XOR2 U1454 ( .A(n1343), .B(n1344), .Z(n1303) );
  ORN2 U1455 ( .A(n1345), .B(n1273), .Z(n1340) );
  AND2 U1456 ( .A(Plaintext[57]), .B(rst), .Z(n1338) );
  ORN2 U1457 ( .A(n1346), .B(n1347), .Z(StateRegInput[56]) );
  AND2 U1458 ( .A(n1348), .B(n1349), .Z(n1347) );
  ORN2 U1459 ( .A(n1249), .B(n1350), .Z(n1349) );
  XOR2 U1460 ( .A(n1311), .B(n1313), .Z(n1350) );
  XOR2 U1461 ( .A(n1351), .B(n1352), .Z(n1311) );
  ORN2 U1462 ( .A(n1353), .B(n1273), .Z(n1348) );
  AND2 U1463 ( .A(Plaintext[56]), .B(rst), .Z(n1346) );
  ORN2 U1464 ( .A(n1354), .B(n1355), .Z(StateRegInput[55]) );
  AND2 U1465 ( .A(n1356), .B(n1357), .Z(n1355) );
  ORN2 U1466 ( .A(n1358), .B(n1261), .Z(n1357) );
  XOR2 U1467 ( .A(n1359), .B(n1327), .Z(n1358) );
  OR2 U1468 ( .A(n1360), .B(n1254), .Z(n1356) );
  AND2 U1469 ( .A(Plaintext[55]), .B(rst), .Z(n1354) );
  ORN2 U1470 ( .A(n1361), .B(n1362), .Z(StateRegInput[54]) );
  AND2 U1471 ( .A(n1363), .B(n1364), .Z(n1362) );
  ORN2 U1472 ( .A(n1249), .B(n1365), .Z(n1364) );
  XOR2 U1473 ( .A(n1366), .B(n1335), .Z(n1365) );
  ORN2 U1474 ( .A(n1254), .B(n1367), .Z(n1363) );
  AND2 U1475 ( .A(Plaintext[54]), .B(rst), .Z(n1361) );
  ORN2 U1476 ( .A(n1368), .B(n1369), .Z(StateRegInput[53]) );
  AND2 U1477 ( .A(n1370), .B(n1371), .Z(n1369) );
  ORN2 U1478 ( .A(n1249), .B(n1372), .Z(n1371) );
  XOR2 U1479 ( .A(n1373), .B(n1344), .Z(n1372) );
  ORN2 U1480 ( .A(n1374), .B(n1273), .Z(n1370) );
  AND2 U1481 ( .A(Plaintext[53]), .B(rst), .Z(n1368) );
  ORN2 U1482 ( .A(n1375), .B(n1376), .Z(StateRegInput[52]) );
  AND2 U1483 ( .A(n1377), .B(n1378), .Z(n1376) );
  ORN2 U1484 ( .A(n1249), .B(n1379), .Z(n1378) );
  XOR2 U1485 ( .A(n1380), .B(n1351), .Z(n1379) );
  ORN2 U1486 ( .A(n1381), .B(n1273), .Z(n1377) );
  AND2 U1487 ( .A(Plaintext[52]), .B(rst), .Z(n1375) );
  ORN2 U1488 ( .A(n1382), .B(n1383), .Z(StateRegInput[51]) );
  AND2 U1489 ( .A(n1384), .B(n1385), .Z(n1383) );
  ORN2 U1490 ( .A(n1249), .B(n1386), .Z(n1385) );
  XOR2 U1491 ( .A(n1359), .B(n1328), .Z(n1386) );
  XOR2 U1492 ( .A(n1289), .B(n1288), .Z(n1359) );
  ORN2 U1493 ( .A(n1387), .B(n1388), .Z(n1289) );
  OR2 U1494 ( .A(n1389), .B(AddKeyConstXOR_XORInst_15_1_N0 ), .Z(n1388) );
  AND2 U1495 ( .A(AddKeyConstXOR_XORInst_15_3_N0 ), .B(
        AddKeyConstXOR_XORInst_15_2_N0 ), .Z(n1389) );
  ORN2 U1496 ( .A(n1254), .B(n1390), .Z(n1384) );
  AND2 U1497 ( .A(Plaintext[51]), .B(rst), .Z(n1382) );
  ORN2 U1498 ( .A(n1391), .B(n1392), .Z(StateRegInput[50]) );
  AND2 U1499 ( .A(n1393), .B(n1394), .Z(n1392) );
  ORN2 U1500 ( .A(n1249), .B(n1395), .Z(n1394) );
  XOR2 U1501 ( .A(n1366), .B(n1336), .Z(n1395) );
  XOR2 U1502 ( .A(n1297), .B(n1296), .Z(n1366) );
  ORN2 U1503 ( .A(n1387), .B(n1396), .Z(n1297) );
  ORN2 U1504 ( .A(n1397), .B(AddKeyConstXOR_XORInst_15_1_N0 ), .Z(n1396) );
  BIC2 U1505 ( .A(n1398), .B(n1399), .Z(n1397) );
  BIC2 U1506 ( .A(n1400), .B(AddKeyConstXOR_XORInst_15_3_N0 ), .Z(n1387) );
  ORN2 U1507 ( .A(n1254), .B(n1401), .Z(n1393) );
  AND2 U1508 ( .A(Plaintext[50]), .B(rst), .Z(n1391) );
  ORN2 U1509 ( .A(n1402), .B(n1403), .Z(StateRegInput[4]) );
  AND2 U1510 ( .A(n1404), .B(n1405), .Z(n1403) );
  ORN2 U1511 ( .A(n1249), .B(n1406), .Z(n1405) );
  XOR2 U1512 ( .A(n1407), .B(n1408), .Z(n1406) );
  ORN2 U1513 ( .A(n1409), .B(n1273), .Z(n1404) );
  AND2 U1514 ( .A(Plaintext[4]), .B(rst), .Z(n1402) );
  ORN2 U1515 ( .A(n1410), .B(n1411), .Z(StateRegInput[49]) );
  AND2 U1516 ( .A(n1412), .B(n1413), .Z(n1411) );
  ORN2 U1517 ( .A(n1414), .B(n1261), .Z(n1413) );
  XOR2 U1518 ( .A(n1373), .B(n1343), .Z(n1414) );
  XOR2 U1519 ( .A(n1304), .B(n1305), .Z(n1373) );
  BIC2 U1520 ( .A(n1415), .B(n1416), .Z(n1305) );
  AND2 U1521 ( .A(n1417), .B(AddKeyConstXOR_XORInst_15_3_N0 ), .Z(n1416) );
  ORN2 U1522 ( .A(n1400), .B(AddKeyConstXOR_XORInst_15_2_N0 ), .Z(n1417) );
  ORN2 U1523 ( .A(AddKeyConstXOR_XORInst_15_0_N1 ), .B(n1398), .Z(n1415) );
  ORN2 U1524 ( .A(n1254), .B(n1418), .Z(n1412) );
  AND2 U1525 ( .A(Plaintext[49]), .B(rst), .Z(n1410) );
  ORN2 U1526 ( .A(n1419), .B(n1420), .Z(StateRegInput[48]) );
  AND2 U1527 ( .A(n1421), .B(n1422), .Z(n1420) );
  ORN2 U1528 ( .A(n1249), .B(n1423), .Z(n1422) );
  XOR2 U1529 ( .A(n1380), .B(n1352), .Z(n1423) );
  XOR2 U1530 ( .A(n1313), .B(n1312), .Z(n1380) );
  ORN2 U1531 ( .A(n1424), .B(n1425), .Z(n1313) );
  AND2 U1532 ( .A(n1426), .B(n1427), .Z(n1425) );
  ORN2 U1533 ( .A(n1398), .B(n1428), .Z(n1427) );
  BIC2 U1534 ( .A(AddKeyConstXOR_XORInst_15_0_N1 ), .B(
        AddKeyConstXOR_XORInst_15_3_N0 ), .Z(n1428) );
  ORN2 U1535 ( .A(AddKeyConstXOR_XORInst_15_2_N0 ), .B(n1399), .Z(n1426) );
  AND2 U1536 ( .A(AddKeyConstXOR_XORInst_15_3_N0 ), .B(
        AddKeyConstXOR_XORInst_15_0_N1 ), .Z(n1399) );
  AND2 U1537 ( .A(AddKeyConstXOR_XORInst_15_1_N0 ), .B(n1429), .Z(n1424) );
  ORN2 U1538 ( .A(n1398), .B(AddKeyConstXOR_XORInst_15_3_N0 ), .Z(n1429) );
  NOT1 U1539 ( .A(AddKeyConstXOR_XORInst_15_2_N0 ), .Z(n1398) );
  ORN2 U1540 ( .A(n1254), .B(n1430), .Z(n1421) );
  AND2 U1541 ( .A(Plaintext[48]), .B(rst), .Z(n1419) );
  ORN2 U1542 ( .A(n1431), .B(n1432), .Z(StateRegInput[47]) );
  AND2 U1543 ( .A(n1433), .B(n1434), .Z(n1432) );
  ORN2 U1544 ( .A(n1435), .B(n1261), .Z(n1434) );
  XOR2 U1545 ( .A(n1436), .B(n1437), .Z(n1435) );
  ORN2 U1546 ( .A(n1437), .B(n1273), .Z(n1433) );
  AND2 U1547 ( .A(Plaintext[47]), .B(rst), .Z(n1431) );
  ORN2 U1548 ( .A(n1438), .B(n1439), .Z(StateRegInput[46]) );
  AND2 U1549 ( .A(n1440), .B(n1441), .Z(n1439) );
  ORN2 U1550 ( .A(n1249), .B(n1442), .Z(n1441) );
  XOR2 U1551 ( .A(n1443), .B(n1444), .Z(n1442) );
  ORN2 U1552 ( .A(n1444), .B(n1273), .Z(n1440) );
  AND2 U1553 ( .A(Plaintext[46]), .B(rst), .Z(n1438) );
  ORN2 U1554 ( .A(n1445), .B(n1446), .Z(StateRegInput[45]) );
  AND2 U1555 ( .A(n1447), .B(n1448), .Z(n1446) );
  ORN2 U1556 ( .A(n1249), .B(n1449), .Z(n1448) );
  XOR2 U1557 ( .A(n1450), .B(n1451), .Z(n1449) );
  OR2 U1558 ( .A(n1451), .B(n1254), .Z(n1447) );
  AND2 U1559 ( .A(Plaintext[45]), .B(rst), .Z(n1445) );
  ORN2 U1560 ( .A(n1452), .B(n1453), .Z(StateRegInput[44]) );
  AND2 U1561 ( .A(n1454), .B(n1455), .Z(n1453) );
  ORN2 U1562 ( .A(n1249), .B(n1456), .Z(n1455) );
  XOR2 U1563 ( .A(n1457), .B(n1458), .Z(n1456) );
  ORN2 U1564 ( .A(n1458), .B(n1273), .Z(n1454) );
  NOT1 U1565 ( .A(n1459), .Z(n1458) );
  AND2 U1566 ( .A(Plaintext[44]), .B(rst), .Z(n1452) );
  ORN2 U1567 ( .A(n1460), .B(n1461), .Z(StateRegInput[43]) );
  AND2 U1568 ( .A(n1462), .B(n1463), .Z(n1461) );
  ORN2 U1569 ( .A(n1464), .B(n1261), .Z(n1463) );
  XOR2 U1570 ( .A(n1436), .B(n1272), .Z(n1464) );
  NOT1 U1571 ( .A(n1465), .Z(n1272) );
  XOR2 U1572 ( .A(n1466), .B(n1467), .Z(n1436) );
  ORN2 U1573 ( .A(n1328), .B(n1273), .Z(n1462) );
  BIC2 U1574 ( .A(n1468), .B(n1469), .Z(n1328) );
  OR2 U1575 ( .A(n1470), .B(AddKeyConstXOR_XORInst_10_1_N0 ), .Z(n1468) );
  AND2 U1576 ( .A(AddKeyConstXOR_XORInst_10_3_N0 ), .B(
        AddKeyConstXOR_XORInst_10_2_N0 ), .Z(n1470) );
  AND2 U1577 ( .A(Plaintext[43]), .B(rst), .Z(n1460) );
  ORN2 U1578 ( .A(n1471), .B(n1472), .Z(StateRegInput[42]) );
  AND2 U1579 ( .A(n1473), .B(n1474), .Z(n1472) );
  ORN2 U1580 ( .A(n1249), .B(n1475), .Z(n1474) );
  XOR2 U1581 ( .A(n1443), .B(n1281), .Z(n1475) );
  NOT1 U1582 ( .A(n1476), .Z(n1281) );
  XOR2 U1583 ( .A(n1477), .B(n1478), .Z(n1443) );
  ORN2 U1584 ( .A(n1336), .B(n1273), .Z(n1473) );
  BIC2 U1585 ( .A(n1479), .B(n1469), .Z(n1336) );
  BIC2 U1586 ( .A(n1480), .B(AddKeyConstXOR_XORInst_10_3_N0 ), .Z(n1469) );
  ORN2 U1587 ( .A(n1481), .B(AddKeyConstXOR_XORInst_10_1_N0 ), .Z(n1479) );
  BIC2 U1588 ( .A(n1482), .B(n1483), .Z(n1481) );
  AND2 U1589 ( .A(Plaintext[42]), .B(rst), .Z(n1471) );
  ORN2 U1590 ( .A(n1484), .B(n1485), .Z(StateRegInput[41]) );
  AND2 U1591 ( .A(n1486), .B(n1487), .Z(n1485) );
  OR2 U1592 ( .A(n1488), .B(n1249), .Z(n1487) );
  XOR2 U1593 ( .A(n1450), .B(n1321), .Z(n1488) );
  XOR2 U1594 ( .A(n1489), .B(n1345), .Z(n1450) );
  ORN2 U1595 ( .A(n1254), .B(n1343), .Z(n1486) );
  BIC2 U1596 ( .A(n1490), .B(n1491), .Z(n1343) );
  AND2 U1597 ( .A(n1492), .B(AddKeyConstXOR_XORInst_10_3_N0 ), .Z(n1491) );
  ORN2 U1598 ( .A(n1480), .B(AddKeyConstXOR_XORInst_10_2_N0 ), .Z(n1492) );
  ORN2 U1599 ( .A(AddKeyConstXOR_XORInst_10_0_N1 ), .B(n1482), .Z(n1490) );
  AND2 U1600 ( .A(Plaintext[41]), .B(rst), .Z(n1484) );
  ORN2 U1601 ( .A(n1493), .B(n1494), .Z(StateRegInput[40]) );
  AND2 U1602 ( .A(n1495), .B(n1496), .Z(n1494) );
  ORN2 U1603 ( .A(n1249), .B(n1497), .Z(n1496) );
  XOR2 U1604 ( .A(n1457), .B(n1409), .Z(n1497) );
  XOR2 U1605 ( .A(n1498), .B(n1499), .Z(n1457) );
  ORN2 U1606 ( .A(n1352), .B(n1273), .Z(n1495) );
  BIC2 U1607 ( .A(n1500), .B(n1501), .Z(n1352) );
  AND2 U1608 ( .A(AddKeyConstXOR_XORInst_10_1_N0 ), .B(n1502), .Z(n1501) );
  ORN2 U1609 ( .A(n1482), .B(AddKeyConstXOR_XORInst_10_3_N0 ), .Z(n1502) );
  AND2 U1610 ( .A(n1503), .B(n1504), .Z(n1500) );
  ORN2 U1611 ( .A(n1482), .B(n1505), .Z(n1504) );
  BIC2 U1612 ( .A(AddKeyConstXOR_XORInst_10_0_N1 ), .B(
        AddKeyConstXOR_XORInst_10_3_N0 ), .Z(n1505) );
  NOT1 U1613 ( .A(AddKeyConstXOR_XORInst_10_2_N0 ), .Z(n1482) );
  ORN2 U1614 ( .A(AddKeyConstXOR_XORInst_10_2_N0 ), .B(n1483), .Z(n1503) );
  AND2 U1615 ( .A(AddKeyConstXOR_XORInst_10_3_N0 ), .B(
        AddKeyConstXOR_XORInst_10_0_N1 ), .Z(n1483) );
  AND2 U1616 ( .A(Plaintext[40]), .B(rst), .Z(n1493) );
  ORN2 U1617 ( .A(n1506), .B(n1507), .Z(StateRegInput[3]) );
  AND2 U1618 ( .A(n1508), .B(n1509), .Z(n1507) );
  ORN2 U1619 ( .A(n1249), .B(n1510), .Z(n1509) );
  XOR2 U1620 ( .A(n1270), .B(n1360), .Z(n1510) );
  XOR2 U1621 ( .A(n1511), .B(n1512), .Z(n1270) );
  ORN2 U1622 ( .A(n1254), .B(n1327), .Z(n1508) );
  BIC2 U1623 ( .A(n1513), .B(n1514), .Z(n1327) );
  AND2 U1624 ( .A(n1515), .B(AddKeyConstXOR_XORInst_0_3_N0 ), .Z(n1514) );
  ORN2 U1625 ( .A(AddKeyConstXOR_XORInst_0_1_N0 ), .B(n1516), .Z(n1515) );
  ORN2 U1626 ( .A(n1517), .B(AddKeyConstXOR_XORInst_0_1_N0 ), .Z(n1513) );
  AND2 U1627 ( .A(Plaintext[3]), .B(rst), .Z(n1506) );
  ORN2 U1628 ( .A(n1518), .B(n1519), .Z(StateRegInput[39]) );
  AND2 U1629 ( .A(n1520), .B(n1521), .Z(n1519) );
  ORN2 U1630 ( .A(n1522), .B(n1261), .Z(n1521) );
  XOR2 U1631 ( .A(n1523), .B(n1329), .Z(n1522) );
  NOT1 U1632 ( .A(n1466), .Z(n1329) );
  ORN2 U1633 ( .A(n1524), .B(n1525), .Z(n1466) );
  ORN2 U1634 ( .A(n1526), .B(AddKeyConstXOR_XORInst_14_1_N0 ), .Z(n1525) );
  AND2 U1635 ( .A(n1527), .B(AddKeyConstXOR_XORInst_14_3_N0 ), .Z(n1524) );
  ORN2 U1636 ( .A(AddKeyConstXOR_XORInst_14_1_N0 ), .B(n1528), .Z(n1527) );
  ORN2 U1637 ( .A(n1529), .B(n1273), .Z(n1520) );
  AND2 U1638 ( .A(Plaintext[39]), .B(rst), .Z(n1518) );
  ORN2 U1639 ( .A(n1530), .B(n1531), .Z(StateRegInput[38]) );
  AND2 U1640 ( .A(n1532), .B(n1533), .Z(n1531) );
  ORN2 U1641 ( .A(n1249), .B(n1534), .Z(n1533) );
  XOR2 U1642 ( .A(n1535), .B(n1337), .Z(n1534) );
  NOT1 U1643 ( .A(n1477), .Z(n1337) );
  ORN2 U1644 ( .A(n1536), .B(n1537), .Z(n1477) );
  ORN2 U1645 ( .A(AddKeyConstXOR_XORInst_14_0_N1 ), .B(n1538), .Z(n1537) );
  AND2 U1646 ( .A(AddKeyConstXOR_XORInst_14_1_N0 ), .B(n1539), .Z(n1536) );
  ORN2 U1647 ( .A(n1540), .B(n1528), .Z(n1539) );
  AND2 U1648 ( .A(AddKeyConstXOR_XORInst_14_3_N0 ), .B(
        AddKeyConstXOR_XORInst_14_0_N1 ), .Z(n1540) );
  ORN2 U1649 ( .A(n1541), .B(n1273), .Z(n1532) );
  AND2 U1650 ( .A(Plaintext[38]), .B(rst), .Z(n1530) );
  ORN2 U1651 ( .A(n1542), .B(n1543), .Z(StateRegInput[37]) );
  AND2 U1652 ( .A(n1544), .B(n1545), .Z(n1543) );
  ORN2 U1653 ( .A(n1249), .B(n1546), .Z(n1545) );
  XOR2 U1654 ( .A(n1547), .B(n1345), .Z(n1546) );
  BIC2 U1655 ( .A(n1548), .B(n1549), .Z(n1345) );
  AND2 U1656 ( .A(n1550), .B(n1538), .Z(n1549) );
  ORN2 U1657 ( .A(AddKeyConstXOR_XORInst_14_0_N1 ), .B(n1528), .Z(n1550) );
  ORN2 U1658 ( .A(n1526), .B(AddKeyConstXOR_XORInst_14_2_N0 ), .Z(n1548) );
  ORN2 U1659 ( .A(n1254), .B(n1551), .Z(n1544) );
  AND2 U1660 ( .A(Plaintext[37]), .B(rst), .Z(n1542) );
  ORN2 U1661 ( .A(n1552), .B(n1553), .Z(StateRegInput[36]) );
  AND2 U1662 ( .A(n1554), .B(n1555), .Z(n1553) );
  ORN2 U1663 ( .A(n1249), .B(n1556), .Z(n1555) );
  XOR2 U1664 ( .A(n1557), .B(n1353), .Z(n1556) );
  NOT1 U1665 ( .A(n1498), .Z(n1353) );
  ORN2 U1666 ( .A(n1558), .B(n1559), .Z(n1498) );
  ORN2 U1667 ( .A(n1560), .B(AddKeyConstXOR_XORInst_14_1_N0 ), .Z(n1559) );
  AND2 U1668 ( .A(AddKeyConstXOR_XORInst_14_2_N0 ), .B(
        AddKeyConstXOR_XORInst_14_3_N0 ), .Z(n1560) );
  AND2 U1669 ( .A(n1561), .B(AddKeyConstXOR_XORInst_14_0_N1 ), .Z(n1558) );
  XOR2 U1670 ( .A(n1528), .B(n1538), .Z(n1561) );
  NOT1 U1671 ( .A(AddKeyConstXOR_XORInst_14_3_N0 ), .Z(n1538) );
  NOT1 U1672 ( .A(AddKeyConstXOR_XORInst_14_2_N0 ), .Z(n1528) );
  ORN2 U1673 ( .A(n1562), .B(n1273), .Z(n1554) );
  AND2 U1674 ( .A(Plaintext[36]), .B(rst), .Z(n1552) );
  ORN2 U1675 ( .A(n1563), .B(n1564), .Z(StateRegInput[35]) );
  AND2 U1676 ( .A(n1565), .B(n1566), .Z(n1564) );
  ORN2 U1677 ( .A(n1249), .B(n1567), .Z(n1566) );
  XOR2 U1678 ( .A(n1523), .B(n1467), .Z(n1567) );
  XOR2 U1679 ( .A(n1465), .B(n1437), .Z(n1523) );
  BIC2 U1680 ( .A(n1568), .B(n1569), .Z(n1437) );
  ORN2 U1681 ( .A(n1570), .B(n1571), .Z(n1568) );
  AND2 U1682 ( .A(AddKeyConstXOR_XORInst_11_3_N0 ), .B(
        AddKeyConstXOR_XORInst_11_2_N0 ), .Z(n1570) );
  ORN2 U1683 ( .A(n1572), .B(n1573), .Z(n1465) );
  OR2 U1684 ( .A(n1574), .B(AddKeyConstXOR_XORInst_1_1_N0 ), .Z(n1573) );
  AND2 U1685 ( .A(AddKeyConstXOR_XORInst_1_3_N0 ), .B(
        AddKeyConstXOR_XORInst_1_2_N0 ), .Z(n1574) );
  ORN2 U1686 ( .A(n1511), .B(n1273), .Z(n1565) );
  AND2 U1687 ( .A(Plaintext[35]), .B(rst), .Z(n1563) );
  ORN2 U1688 ( .A(n1575), .B(n1576), .Z(StateRegInput[34]) );
  AND2 U1689 ( .A(n1577), .B(n1578), .Z(n1576) );
  ORN2 U1690 ( .A(n1249), .B(n1579), .Z(n1578) );
  XOR2 U1691 ( .A(n1535), .B(n1478), .Z(n1579) );
  XOR2 U1692 ( .A(n1476), .B(n1444), .Z(n1535) );
  BIC2 U1693 ( .A(n1580), .B(n1569), .Z(n1444) );
  BIC2 U1694 ( .A(n1581), .B(AddKeyConstXOR_XORInst_11_3_N0 ), .Z(n1569) );
  ORN2 U1695 ( .A(n1582), .B(AddKeyConstXOR_XORInst_11_1_N0 ), .Z(n1580) );
  BIC2 U1696 ( .A(n1583), .B(n1584), .Z(n1582) );
  ORN2 U1697 ( .A(n1572), .B(n1585), .Z(n1476) );
  ORN2 U1698 ( .A(n1586), .B(AddKeyConstXOR_XORInst_1_1_N0 ), .Z(n1585) );
  BIC2 U1699 ( .A(n1587), .B(n1588), .Z(n1586) );
  BIC2 U1700 ( .A(n1589), .B(AddKeyConstXOR_XORInst_1_3_N0 ), .Z(n1572) );
  ORN2 U1701 ( .A(n1590), .B(n1273), .Z(n1577) );
  AND2 U1702 ( .A(Plaintext[34]), .B(rst), .Z(n1575) );
  ORN2 U1703 ( .A(n1591), .B(n1592), .Z(StateRegInput[33]) );
  AND2 U1704 ( .A(n1593), .B(n1594), .Z(n1592) );
  ORN2 U1705 ( .A(n1595), .B(n1261), .Z(n1594) );
  XOR2 U1706 ( .A(n1547), .B(n1489), .Z(n1595) );
  XOR2 U1707 ( .A(n1451), .B(n1321), .Z(n1547) );
  BIC2 U1708 ( .A(n1596), .B(n1597), .Z(n1321) );
  AND2 U1709 ( .A(n1598), .B(AddKeyConstXOR_XORInst_1_3_N0 ), .Z(n1597) );
  ORN2 U1710 ( .A(n1589), .B(AddKeyConstXOR_XORInst_1_2_N0 ), .Z(n1598) );
  ORN2 U1711 ( .A(AddKeyConstXOR_XORInst_1_0_N1 ), .B(n1587), .Z(n1596) );
  ORN2 U1712 ( .A(n1599), .B(n1600), .Z(n1451) );
  ORN2 U1713 ( .A(AddKeyConstXOR_XORInst_11_0_N1 ), .B(n1583), .Z(n1600) );
  AND2 U1714 ( .A(n1601), .B(AddKeyConstXOR_XORInst_11_3_N0 ), .Z(n1599) );
  ORN2 U1715 ( .A(n1253), .B(n1273), .Z(n1593) );
  AND2 U1716 ( .A(Plaintext[33]), .B(rst), .Z(n1591) );
  ORN2 U1717 ( .A(n1602), .B(n1603), .Z(StateRegInput[32]) );
  AND2 U1718 ( .A(n1604), .B(n1605), .Z(n1603) );
  ORN2 U1719 ( .A(n1249), .B(n1606), .Z(n1605) );
  XOR2 U1720 ( .A(n1557), .B(n1499), .Z(n1606) );
  XOR2 U1721 ( .A(n1459), .B(n1409), .Z(n1557) );
  BIC2 U1722 ( .A(n1607), .B(n1608), .Z(n1409) );
  AND2 U1723 ( .A(AddKeyConstXOR_XORInst_1_1_N0 ), .B(n1609), .Z(n1608) );
  ORN2 U1724 ( .A(n1587), .B(AddKeyConstXOR_XORInst_1_3_N0 ), .Z(n1609) );
  AND2 U1725 ( .A(n1610), .B(n1611), .Z(n1607) );
  ORN2 U1726 ( .A(n1587), .B(n1612), .Z(n1611) );
  BIC2 U1727 ( .A(AddKeyConstXOR_XORInst_1_0_N1 ), .B(
        AddKeyConstXOR_XORInst_1_3_N0 ), .Z(n1612) );
  NOT1 U1728 ( .A(AddKeyConstXOR_XORInst_1_2_N0 ), .Z(n1587) );
  ORN2 U1729 ( .A(AddKeyConstXOR_XORInst_1_2_N0 ), .B(n1588), .Z(n1610) );
  AND2 U1730 ( .A(AddKeyConstXOR_XORInst_1_3_N0 ), .B(
        AddKeyConstXOR_XORInst_1_0_N1 ), .Z(n1588) );
  ORN2 U1731 ( .A(n1613), .B(n1614), .Z(n1459) );
  OR2 U1732 ( .A(n1615), .B(AddKeyConstXOR_XORInst_11_3_N0 ), .Z(n1614) );
  AND2 U1733 ( .A(n1601), .B(n1571), .Z(n1615) );
  ORN2 U1734 ( .A(n1581), .B(AddKeyConstXOR_XORInst_11_2_N0 ), .Z(n1601) );
  AND2 U1735 ( .A(n1616), .B(n1583), .Z(n1613) );
  NOT1 U1736 ( .A(AddKeyConstXOR_XORInst_11_2_N0 ), .Z(n1583) );
  ORN2 U1737 ( .A(n1584), .B(n1571), .Z(n1616) );
  NOT1 U1738 ( .A(AddKeyConstXOR_XORInst_11_1_N0 ), .Z(n1571) );
  AND2 U1739 ( .A(AddKeyConstXOR_XORInst_11_3_N0 ), .B(
        AddKeyConstXOR_XORInst_11_0_N1 ), .Z(n1584) );
  ORN2 U1740 ( .A(n1263), .B(n1273), .Z(n1604) );
  AND2 U1741 ( .A(Plaintext[32]), .B(rst), .Z(n1602) );
  ORN2 U1742 ( .A(n1617), .B(n1618), .Z(StateRegInput[31]) );
  AND2 U1743 ( .A(n1619), .B(n1620), .Z(n1618) );
  ORN2 U1744 ( .A(n1621), .B(n1261), .Z(n1620) );
  XOR2 U1745 ( .A(n1622), .B(n1390), .Z(n1621) );
  ORN2 U1746 ( .A(n1254), .B(n1271), .Z(n1619) );
  AND2 U1747 ( .A(Plaintext[31]), .B(rst), .Z(n1617) );
  ORN2 U1748 ( .A(n1623), .B(n1624), .Z(StateRegInput[30]) );
  AND2 U1749 ( .A(n1625), .B(n1626), .Z(n1624) );
  ORN2 U1750 ( .A(n1249), .B(n1627), .Z(n1626) );
  XOR2 U1751 ( .A(n1628), .B(n1401), .Z(n1627) );
  ORN2 U1752 ( .A(n1280), .B(n1273), .Z(n1625) );
  AND2 U1753 ( .A(Plaintext[30]), .B(rst), .Z(n1623) );
  ORN2 U1754 ( .A(n1629), .B(n1630), .Z(StateRegInput[2]) );
  AND2 U1755 ( .A(n1631), .B(n1632), .Z(n1630) );
  ORN2 U1756 ( .A(n1249), .B(n1633), .Z(n1632) );
  XOR2 U1757 ( .A(n1279), .B(n1367), .Z(n1633) );
  XOR2 U1758 ( .A(n1590), .B(n1634), .Z(n1279) );
  ORN2 U1759 ( .A(n1335), .B(n1273), .Z(n1631) );
  BIC2 U1760 ( .A(n1635), .B(n1636), .Z(n1335) );
  AND2 U1761 ( .A(n1637), .B(AddKeyConstXOR_XORInst_0_1_N0 ), .Z(n1636) );
  ORN2 U1762 ( .A(n1638), .B(n1516), .Z(n1637) );
  OR2 U1763 ( .A(AddKeyConstXOR_XORInst_0_3_N0 ), .B(
        AddKeyConstXOR_XORInst_0_0_N1 ), .Z(n1635) );
  AND2 U1764 ( .A(Plaintext[2]), .B(rst), .Z(n1629) );
  ORN2 U1765 ( .A(n1639), .B(n1640), .Z(StateRegInput[29]) );
  AND2 U1766 ( .A(n1641), .B(n1642), .Z(n1640) );
  ORN2 U1767 ( .A(n1643), .B(n1261), .Z(n1642) );
  XOR2 U1768 ( .A(n1644), .B(n1418), .Z(n1643) );
  ORN2 U1769 ( .A(n1320), .B(n1273), .Z(n1641) );
  AND2 U1770 ( .A(Plaintext[29]), .B(rst), .Z(n1639) );
  ORN2 U1771 ( .A(n1645), .B(n1646), .Z(StateRegInput[28]) );
  AND2 U1772 ( .A(n1647), .B(n1648), .Z(n1646) );
  ORN2 U1773 ( .A(n1249), .B(n1649), .Z(n1648) );
  XOR2 U1774 ( .A(n1650), .B(n1430), .Z(n1649) );
  ORN2 U1775 ( .A(n1408), .B(n1273), .Z(n1647) );
  AND2 U1776 ( .A(Plaintext[28]), .B(rst), .Z(n1645) );
  ORN2 U1777 ( .A(n1651), .B(n1652), .Z(StateRegInput[27]) );
  AND2 U1778 ( .A(n1653), .B(n1654), .Z(n1652) );
  ORN2 U1779 ( .A(n1249), .B(n1655), .Z(n1654) );
  XOR2 U1780 ( .A(n1622), .B(n1656), .Z(n1655) );
  XOR2 U1781 ( .A(n1657), .B(n1529), .Z(n1622) );
  ORN2 U1782 ( .A(n1656), .B(n1273), .Z(n1653) );
  AND2 U1783 ( .A(Plaintext[27]), .B(rst), .Z(n1651) );
  ORN2 U1784 ( .A(n1658), .B(n1659), .Z(StateRegInput[26]) );
  AND2 U1785 ( .A(n1660), .B(n1661), .Z(n1659) );
  OR2 U1786 ( .A(n1662), .B(n1249), .Z(n1661) );
  XOR2 U1787 ( .A(n1628), .B(n1663), .Z(n1662) );
  XOR2 U1788 ( .A(n1664), .B(n1541), .Z(n1628) );
  ORN2 U1789 ( .A(n1663), .B(n1273), .Z(n1660) );
  AND2 U1790 ( .A(Plaintext[26]), .B(rst), .Z(n1658) );
  ORN2 U1791 ( .A(n1665), .B(n1666), .Z(StateRegInput[25]) );
  AND2 U1792 ( .A(n1667), .B(n1668), .Z(n1666) );
  ORN2 U1793 ( .A(n1249), .B(n1669), .Z(n1668) );
  XOR2 U1794 ( .A(n1644), .B(n1670), .Z(n1669) );
  XOR2 U1795 ( .A(n1671), .B(n1551), .Z(n1644) );
  OR2 U1796 ( .A(n1670), .B(n1254), .Z(n1667) );
  AND2 U1797 ( .A(Plaintext[25]), .B(rst), .Z(n1665) );
  ORN2 U1798 ( .A(n1672), .B(n1673), .Z(StateRegInput[24]) );
  AND2 U1799 ( .A(n1674), .B(n1675), .Z(n1673) );
  OR2 U1800 ( .A(n1676), .B(n1249), .Z(n1675) );
  XOR2 U1801 ( .A(n1650), .B(n1677), .Z(n1676) );
  XOR2 U1802 ( .A(n1678), .B(n1562), .Z(n1650) );
  ORN2 U1803 ( .A(n1677), .B(n1273), .Z(n1674) );
  AND2 U1804 ( .A(Plaintext[24]), .B(rst), .Z(n1672) );
  ORN2 U1805 ( .A(n1679), .B(n1680), .Z(StateRegInput[23]) );
  AND2 U1806 ( .A(n1681), .B(n1682), .Z(n1680) );
  ORN2 U1807 ( .A(n1249), .B(n1683), .Z(n1682) );
  XOR2 U1808 ( .A(n1684), .B(n1529), .Z(n1683) );
  BIC2 U1809 ( .A(n1685), .B(n1686), .Z(n1529) );
  OR2 U1810 ( .A(n1687), .B(AddKeyConstXOR_XORInst_9_1_N0 ), .Z(n1685) );
  AND2 U1811 ( .A(AddKeyConstXOR_XORInst_9_3_N0 ), .B(
        AddKeyConstXOR_XORInst_9_2_N0 ), .Z(n1687) );
  ORN2 U1812 ( .A(n1288), .B(n1273), .Z(n1681) );
  BIC2 U1813 ( .A(n1688), .B(n1689), .Z(n1288) );
  OR2 U1814 ( .A(n1690), .B(AddKeyConstXOR_XORInst_5_1_N0 ), .Z(n1688) );
  AND2 U1815 ( .A(AddKeyConstXOR_XORInst_5_3_N0 ), .B(
        AddKeyConstXOR_XORInst_5_2_N0 ), .Z(n1690) );
  AND2 U1816 ( .A(Plaintext[23]), .B(rst), .Z(n1679) );
  ORN2 U1817 ( .A(n1691), .B(n1692), .Z(StateRegInput[22]) );
  AND2 U1818 ( .A(n1693), .B(n1694), .Z(n1692) );
  ORN2 U1819 ( .A(n1249), .B(n1695), .Z(n1694) );
  XOR2 U1820 ( .A(n1696), .B(n1541), .Z(n1695) );
  BIC2 U1821 ( .A(n1697), .B(n1686), .Z(n1541) );
  BIC2 U1822 ( .A(n1698), .B(AddKeyConstXOR_XORInst_9_3_N0 ), .Z(n1686) );
  ORN2 U1823 ( .A(n1699), .B(AddKeyConstXOR_XORInst_9_1_N0 ), .Z(n1697) );
  BIC2 U1824 ( .A(n1700), .B(n1701), .Z(n1699) );
  ORN2 U1825 ( .A(n1296), .B(n1273), .Z(n1693) );
  BIC2 U1826 ( .A(n1702), .B(n1689), .Z(n1296) );
  BIC2 U1827 ( .A(n1703), .B(AddKeyConstXOR_XORInst_5_3_N0 ), .Z(n1689) );
  ORN2 U1828 ( .A(n1704), .B(AddKeyConstXOR_XORInst_5_1_N0 ), .Z(n1702) );
  BIC2 U1829 ( .A(n1705), .B(n1706), .Z(n1704) );
  AND2 U1830 ( .A(Plaintext[22]), .B(rst), .Z(n1691) );
  ORN2 U1831 ( .A(n1707), .B(n1708), .Z(StateRegInput[21]) );
  AND2 U1832 ( .A(n1709), .B(n1710), .Z(n1708) );
  ORN2 U1833 ( .A(n1711), .B(n1261), .Z(n1710) );
  XOR2 U1834 ( .A(n1712), .B(n1551), .Z(n1711) );
  BIC2 U1835 ( .A(n1713), .B(n1714), .Z(n1551) );
  AND2 U1836 ( .A(n1715), .B(AddKeyConstXOR_XORInst_9_3_N0 ), .Z(n1714) );
  ORN2 U1837 ( .A(n1698), .B(AddKeyConstXOR_XORInst_9_2_N0 ), .Z(n1715) );
  ORN2 U1838 ( .A(AddKeyConstXOR_XORInst_9_0_N1 ), .B(n1700), .Z(n1713) );
  OR2 U1839 ( .A(n1304), .B(n1254), .Z(n1709) );
  ORN2 U1840 ( .A(n1716), .B(n1717), .Z(n1304) );
  ORN2 U1841 ( .A(AddKeyConstXOR_XORInst_5_0_N1 ), .B(n1705), .Z(n1717) );
  AND2 U1842 ( .A(n1718), .B(AddKeyConstXOR_XORInst_5_3_N0 ), .Z(n1716) );
  ORN2 U1843 ( .A(n1703), .B(AddKeyConstXOR_XORInst_5_2_N0 ), .Z(n1718) );
  AND2 U1844 ( .A(Plaintext[21]), .B(rst), .Z(n1707) );
  ORN2 U1845 ( .A(n1719), .B(n1720), .Z(StateRegInput[20]) );
  AND2 U1846 ( .A(n1721), .B(n1722), .Z(n1720) );
  ORN2 U1847 ( .A(n1249), .B(n1723), .Z(n1722) );
  XOR2 U1848 ( .A(n1724), .B(n1562), .Z(n1723) );
  BIC2 U1849 ( .A(n1725), .B(n1726), .Z(n1562) );
  AND2 U1850 ( .A(AddKeyConstXOR_XORInst_9_1_N0 ), .B(n1727), .Z(n1726) );
  ORN2 U1851 ( .A(n1700), .B(AddKeyConstXOR_XORInst_9_3_N0 ), .Z(n1727) );
  AND2 U1852 ( .A(n1728), .B(n1729), .Z(n1725) );
  ORN2 U1853 ( .A(n1700), .B(n1730), .Z(n1729) );
  BIC2 U1854 ( .A(AddKeyConstXOR_XORInst_9_0_N1 ), .B(
        AddKeyConstXOR_XORInst_9_3_N0 ), .Z(n1730) );
  NOT1 U1855 ( .A(AddKeyConstXOR_XORInst_9_2_N0 ), .Z(n1700) );
  ORN2 U1856 ( .A(AddKeyConstXOR_XORInst_9_2_N0 ), .B(n1701), .Z(n1728) );
  AND2 U1857 ( .A(AddKeyConstXOR_XORInst_9_3_N0 ), .B(
        AddKeyConstXOR_XORInst_9_0_N1 ), .Z(n1701) );
  ORN2 U1858 ( .A(n1312), .B(n1273), .Z(n1721) );
  BIC2 U1859 ( .A(n1731), .B(n1732), .Z(n1312) );
  AND2 U1860 ( .A(AddKeyConstXOR_XORInst_5_1_N0 ), .B(n1733), .Z(n1732) );
  ORN2 U1861 ( .A(n1705), .B(AddKeyConstXOR_XORInst_5_3_N0 ), .Z(n1733) );
  AND2 U1862 ( .A(n1734), .B(n1735), .Z(n1731) );
  ORN2 U1863 ( .A(n1705), .B(n1736), .Z(n1735) );
  BIC2 U1864 ( .A(AddKeyConstXOR_XORInst_5_0_N1 ), .B(
        AddKeyConstXOR_XORInst_5_3_N0 ), .Z(n1736) );
  NOT1 U1865 ( .A(AddKeyConstXOR_XORInst_5_2_N0 ), .Z(n1705) );
  ORN2 U1866 ( .A(AddKeyConstXOR_XORInst_5_2_N0 ), .B(n1706), .Z(n1734) );
  AND2 U1867 ( .A(AddKeyConstXOR_XORInst_5_3_N0 ), .B(
        AddKeyConstXOR_XORInst_5_0_N1 ), .Z(n1706) );
  AND2 U1868 ( .A(Plaintext[20]), .B(rst), .Z(n1719) );
  ORN2 U1869 ( .A(n1737), .B(n1738), .Z(StateRegInput[1]) );
  AND2 U1870 ( .A(n1739), .B(n1740), .Z(n1738) );
  ORN2 U1871 ( .A(n1249), .B(n1741), .Z(n1740) );
  XOR2 U1872 ( .A(n1319), .B(n1374), .Z(n1741) );
  XOR2 U1873 ( .A(n1253), .B(n1255), .Z(n1319) );
  ORN2 U1874 ( .A(n1742), .B(n1743), .Z(n1253) );
  ORN2 U1875 ( .A(AddKeyConstXOR_XORInst_8_0_N1 ), .B(n1744), .Z(n1743) );
  AND2 U1876 ( .A(n1745), .B(AddKeyConstXOR_XORInst_8_3_N0 ), .Z(n1742) );
  ORN2 U1877 ( .A(n1746), .B(AddKeyConstXOR_XORInst_8_2_N0 ), .Z(n1745) );
  ORN2 U1878 ( .A(n1344), .B(n1273), .Z(n1739) );
  BIC2 U1879 ( .A(n1747), .B(n1748), .Z(n1344) );
  BIC2 U1880 ( .A(n1749), .B(AddKeyConstXOR_XORInst_0_3_N0 ), .Z(n1748) );
  ORN2 U1881 ( .A(AddKeyConstXOR_XORInst_0_0_N1 ), .B(n1516), .Z(n1749) );
  AND2 U1882 ( .A(Plaintext[1]), .B(rst), .Z(n1737) );
  ORN2 U1883 ( .A(n1750), .B(n1751), .Z(StateRegInput[19]) );
  AND2 U1884 ( .A(n1752), .B(n1753), .Z(n1751) );
  ORN2 U1885 ( .A(n1754), .B(n1261), .Z(n1753) );
  XOR2 U1886 ( .A(n1684), .B(n1657), .Z(n1754) );
  XOR2 U1887 ( .A(n1390), .B(n1656), .Z(n1684) );
  BIC2 U1888 ( .A(n1755), .B(n1756), .Z(n1656) );
  OR2 U1889 ( .A(n1757), .B(AddKeyConstXOR_XORInst_6_1_N0 ), .Z(n1755) );
  AND2 U1890 ( .A(AddKeyConstXOR_XORInst_6_3_N0 ), .B(
        AddKeyConstXOR_XORInst_6_2_N0 ), .Z(n1757) );
  ORN2 U1891 ( .A(n1758), .B(n1759), .Z(n1390) );
  OR2 U1892 ( .A(n1760), .B(AddKeyConstXOR_XORInst_12_1_N0 ), .Z(n1759) );
  AND2 U1893 ( .A(AddKeyConstXOR_XORInst_12_3_N0 ), .B(
        AddKeyConstXOR_XORInst_12_2_N0 ), .Z(n1760) );
  ORN2 U1894 ( .A(n1467), .B(n1273), .Z(n1752) );
  BIC2 U1895 ( .A(n1761), .B(n1762), .Z(n1467) );
  OR2 U1896 ( .A(n1763), .B(AddKeyConstXOR_XORInst_4_1_N0 ), .Z(n1761) );
  AND2 U1897 ( .A(AddKeyConstXOR_XORInst_4_3_N0 ), .B(
        AddKeyConstXOR_XORInst_4_2_N0 ), .Z(n1763) );
  AND2 U1898 ( .A(Plaintext[19]), .B(rst), .Z(n1750) );
  ORN2 U1899 ( .A(n1764), .B(n1765), .Z(StateRegInput[18]) );
  AND2 U1900 ( .A(n1766), .B(n1767), .Z(n1765) );
  ORN2 U1901 ( .A(n1249), .B(n1768), .Z(n1767) );
  XOR2 U1902 ( .A(n1696), .B(n1664), .Z(n1768) );
  XOR2 U1903 ( .A(n1401), .B(n1663), .Z(n1696) );
  BIC2 U1904 ( .A(n1769), .B(n1756), .Z(n1663) );
  BIC2 U1905 ( .A(n1770), .B(AddKeyConstXOR_XORInst_6_3_N0 ), .Z(n1756) );
  ORN2 U1906 ( .A(n1771), .B(AddKeyConstXOR_XORInst_6_1_N0 ), .Z(n1769) );
  BIC2 U1907 ( .A(n1772), .B(n1773), .Z(n1771) );
  ORN2 U1908 ( .A(n1758), .B(n1774), .Z(n1401) );
  ORN2 U1909 ( .A(n1775), .B(AddKeyConstXOR_XORInst_12_1_N0 ), .Z(n1774) );
  BIC2 U1910 ( .A(n1776), .B(n1777), .Z(n1775) );
  BIC2 U1911 ( .A(n1778), .B(AddKeyConstXOR_XORInst_12_3_N0 ), .Z(n1758) );
  ORN2 U1912 ( .A(n1478), .B(n1273), .Z(n1766) );
  BIC2 U1913 ( .A(n1779), .B(n1762), .Z(n1478) );
  BIC2 U1914 ( .A(n1780), .B(AddKeyConstXOR_XORInst_4_3_N0 ), .Z(n1762) );
  ORN2 U1915 ( .A(n1781), .B(AddKeyConstXOR_XORInst_4_1_N0 ), .Z(n1779) );
  BIC2 U1916 ( .A(n1782), .B(n1783), .Z(n1781) );
  AND2 U1917 ( .A(Plaintext[18]), .B(rst), .Z(n1764) );
  ORN2 U1918 ( .A(n1784), .B(n1785), .Z(StateRegInput[17]) );
  AND2 U1919 ( .A(n1786), .B(n1787), .Z(n1785) );
  ORN2 U1920 ( .A(n1249), .B(n1788), .Z(n1787) );
  XOR2 U1921 ( .A(n1712), .B(n1671), .Z(n1788) );
  XOR2 U1922 ( .A(n1670), .B(n1418), .Z(n1712) );
  BIC2 U1923 ( .A(n1789), .B(n1790), .Z(n1418) );
  AND2 U1924 ( .A(n1791), .B(AddKeyConstXOR_XORInst_12_3_N0 ), .Z(n1790) );
  ORN2 U1925 ( .A(n1778), .B(AddKeyConstXOR_XORInst_12_2_N0 ), .Z(n1791) );
  ORN2 U1926 ( .A(AddKeyConstXOR_XORInst_12_0_N1 ), .B(n1776), .Z(n1789) );
  ORN2 U1927 ( .A(n1792), .B(n1793), .Z(n1670) );
  ORN2 U1928 ( .A(AddKeyConstXOR_XORInst_6_0_N1 ), .B(n1772), .Z(n1793) );
  AND2 U1929 ( .A(n1794), .B(AddKeyConstXOR_XORInst_6_3_N0 ), .Z(n1792) );
  ORN2 U1930 ( .A(n1770), .B(AddKeyConstXOR_XORInst_6_2_N0 ), .Z(n1794) );
  ORN2 U1931 ( .A(n1254), .B(n1489), .Z(n1786) );
  BIC2 U1932 ( .A(n1795), .B(n1796), .Z(n1489) );
  AND2 U1933 ( .A(n1797), .B(AddKeyConstXOR_XORInst_4_3_N0 ), .Z(n1796) );
  ORN2 U1934 ( .A(n1780), .B(AddKeyConstXOR_XORInst_4_2_N0 ), .Z(n1797) );
  ORN2 U1935 ( .A(AddKeyConstXOR_XORInst_4_0_N1 ), .B(n1782), .Z(n1795) );
  AND2 U1936 ( .A(Plaintext[17]), .B(rst), .Z(n1784) );
  ORN2 U1937 ( .A(n1798), .B(n1799), .Z(StateRegInput[16]) );
  AND2 U1938 ( .A(n1800), .B(n1801), .Z(n1799) );
  ORN2 U1939 ( .A(n1249), .B(n1802), .Z(n1801) );
  XOR2 U1940 ( .A(n1724), .B(n1678), .Z(n1802) );
  XOR2 U1941 ( .A(n1430), .B(n1677), .Z(n1724) );
  BIC2 U1942 ( .A(n1803), .B(n1804), .Z(n1677) );
  AND2 U1943 ( .A(AddKeyConstXOR_XORInst_6_1_N0 ), .B(n1805), .Z(n1804) );
  ORN2 U1944 ( .A(n1772), .B(AddKeyConstXOR_XORInst_6_3_N0 ), .Z(n1805) );
  AND2 U1945 ( .A(n1806), .B(n1807), .Z(n1803) );
  ORN2 U1946 ( .A(n1772), .B(n1808), .Z(n1807) );
  BIC2 U1947 ( .A(AddKeyConstXOR_XORInst_6_0_N1 ), .B(
        AddKeyConstXOR_XORInst_6_3_N0 ), .Z(n1808) );
  NOT1 U1948 ( .A(AddKeyConstXOR_XORInst_6_2_N0 ), .Z(n1772) );
  ORN2 U1949 ( .A(AddKeyConstXOR_XORInst_6_2_N0 ), .B(n1773), .Z(n1806) );
  AND2 U1950 ( .A(AddKeyConstXOR_XORInst_6_3_N0 ), .B(
        AddKeyConstXOR_XORInst_6_0_N1 ), .Z(n1773) );
  ORN2 U1951 ( .A(n1809), .B(n1810), .Z(n1430) );
  AND2 U1952 ( .A(n1811), .B(n1812), .Z(n1810) );
  ORN2 U1953 ( .A(n1776), .B(n1813), .Z(n1812) );
  BIC2 U1954 ( .A(AddKeyConstXOR_XORInst_12_0_N1 ), .B(
        AddKeyConstXOR_XORInst_12_3_N0 ), .Z(n1813) );
  ORN2 U1955 ( .A(AddKeyConstXOR_XORInst_12_2_N0 ), .B(n1777), .Z(n1811) );
  AND2 U1956 ( .A(AddKeyConstXOR_XORInst_12_3_N0 ), .B(
        AddKeyConstXOR_XORInst_12_0_N1 ), .Z(n1777) );
  AND2 U1957 ( .A(AddKeyConstXOR_XORInst_12_1_N0 ), .B(n1814), .Z(n1809) );
  ORN2 U1958 ( .A(n1776), .B(AddKeyConstXOR_XORInst_12_3_N0 ), .Z(n1814) );
  NOT1 U1959 ( .A(AddKeyConstXOR_XORInst_12_2_N0 ), .Z(n1776) );
  ORN2 U1960 ( .A(n1499), .B(n1273), .Z(n1800) );
  BIC2 U1961 ( .A(n1815), .B(n1816), .Z(n1499) );
  AND2 U1962 ( .A(AddKeyConstXOR_XORInst_4_1_N0 ), .B(n1817), .Z(n1816) );
  ORN2 U1963 ( .A(n1782), .B(AddKeyConstXOR_XORInst_4_3_N0 ), .Z(n1817) );
  AND2 U1964 ( .A(n1818), .B(n1819), .Z(n1815) );
  ORN2 U1965 ( .A(n1782), .B(n1820), .Z(n1819) );
  BIC2 U1966 ( .A(AddKeyConstXOR_XORInst_4_0_N1 ), .B(
        AddKeyConstXOR_XORInst_4_3_N0 ), .Z(n1820) );
  NOT1 U1967 ( .A(AddKeyConstXOR_XORInst_4_2_N0 ), .Z(n1782) );
  ORN2 U1968 ( .A(AddKeyConstXOR_XORInst_4_2_N0 ), .B(n1783), .Z(n1818) );
  AND2 U1969 ( .A(AddKeyConstXOR_XORInst_4_3_N0 ), .B(
        AddKeyConstXOR_XORInst_4_0_N1 ), .Z(n1783) );
  AND2 U1970 ( .A(Plaintext[16]), .B(rst), .Z(n1798) );
  ORN2 U1971 ( .A(n1821), .B(n1822), .Z(StateRegInput[15]) );
  AND2 U1972 ( .A(n1823), .B(n1824), .Z(n1822) );
  ORN2 U1973 ( .A(n1825), .B(n1261), .Z(n1824) );
  NOT1 U1974 ( .A(n1249), .Z(n1261) );
  XOR2 U1975 ( .A(n1826), .B(n1512), .Z(n1825) );
  ORN2 U1976 ( .A(n1254), .B(n1657), .Z(n1823) );
  BIC2 U1977 ( .A(n1827), .B(n1828), .Z(n1657) );
  AND2 U1978 ( .A(n1829), .B(AddKeyConstXOR_XORInst_3_3_N0 ), .Z(n1828) );
  ORN2 U1979 ( .A(AddKeyConstXOR_XORInst_3_1_N0 ), .B(n1830), .Z(n1829) );
  ORN2 U1980 ( .A(n1831), .B(AddKeyConstXOR_XORInst_3_1_N0 ), .Z(n1827) );
  AND2 U1981 ( .A(Plaintext[15]), .B(rst), .Z(n1821) );
  ORN2 U1982 ( .A(n1832), .B(n1833), .Z(StateRegInput[14]) );
  AND2 U1983 ( .A(n1834), .B(n1835), .Z(n1833) );
  ORN2 U1984 ( .A(n1249), .B(n1836), .Z(n1835) );
  XOR2 U1985 ( .A(n1837), .B(n1634), .Z(n1836) );
  ORN2 U1986 ( .A(n1664), .B(n1273), .Z(n1834) );
  BIC2 U1987 ( .A(n1838), .B(n1839), .Z(n1664) );
  AND2 U1988 ( .A(n1840), .B(AddKeyConstXOR_XORInst_3_1_N0 ), .Z(n1839) );
  ORN2 U1989 ( .A(n1841), .B(n1830), .Z(n1840) );
  OR2 U1990 ( .A(AddKeyConstXOR_XORInst_3_3_N0 ), .B(
        AddKeyConstXOR_XORInst_3_0_N1 ), .Z(n1838) );
  AND2 U1991 ( .A(Plaintext[14]), .B(rst), .Z(n1832) );
  ORN2 U1992 ( .A(n1842), .B(n1843), .Z(StateRegInput[13]) );
  AND2 U1993 ( .A(n1844), .B(n1845), .Z(n1843) );
  ORN2 U1994 ( .A(n1249), .B(n1846), .Z(n1845) );
  XOR2 U1995 ( .A(n1251), .B(n1255), .Z(n1846) );
  BIC2 U1996 ( .A(n1847), .B(n1848), .Z(n1255) );
  AND2 U1997 ( .A(n1849), .B(AddKeyConstXOR_XORInst_2_3_N0 ), .Z(n1848) );
  ORN2 U1998 ( .A(n1850), .B(AddKeyConstXOR_XORInst_2_2_N0 ), .Z(n1849) );
  ORN2 U1999 ( .A(AddKeyConstXOR_XORInst_2_0_N1 ), .B(n1851), .Z(n1847) );
  XOR2 U2000 ( .A(n1374), .B(n1320), .Z(n1251) );
  BIC2 U2001 ( .A(n1852), .B(n1853), .Z(n1320) );
  BIC2 U2002 ( .A(n1854), .B(AddKeyConstXOR_XORInst_7_3_N0 ), .Z(n1853) );
  ORN2 U2003 ( .A(AddKeyConstXOR_XORInst_7_0_N1 ), .B(n1855), .Z(n1854) );
  ORN2 U2004 ( .A(n1856), .B(n1857), .Z(n1374) );
  ORN2 U2005 ( .A(AddKeyConstXOR_XORInst_13_0_N1 ), .B(n1858), .Z(n1857) );
  AND2 U2006 ( .A(n1859), .B(AddKeyConstXOR_XORInst_13_3_N0 ), .Z(n1856) );
  ORN2 U2007 ( .A(n1860), .B(AddKeyConstXOR_XORInst_13_2_N0 ), .Z(n1859) );
  ORN2 U2008 ( .A(n1671), .B(n1273), .Z(n1844) );
  BIC2 U2009 ( .A(n1861), .B(n1862), .Z(n1671) );
  BIC2 U2010 ( .A(n1863), .B(AddKeyConstXOR_XORInst_3_3_N0 ), .Z(n1862) );
  ORN2 U2011 ( .A(AddKeyConstXOR_XORInst_3_0_N1 ), .B(n1830), .Z(n1863) );
  AND2 U2012 ( .A(Plaintext[13]), .B(rst), .Z(n1842) );
  ORN2 U2013 ( .A(n1864), .B(n1865), .Z(StateRegInput[12]) );
  AND2 U2014 ( .A(n1866), .B(n1867), .Z(n1865) );
  ORN2 U2015 ( .A(n1249), .B(n1868), .Z(n1867) );
  XOR2 U2016 ( .A(n1262), .B(n1264), .Z(n1868) );
  XOR2 U2017 ( .A(n1408), .B(n1381), .Z(n1262) );
  BIC2 U2018 ( .A(n1869), .B(n1870), .Z(n1408) );
  AND2 U2019 ( .A(n1871), .B(n1855), .Z(n1870) );
  OR2 U2020 ( .A(n1872), .B(AddKeyConstXOR_XORInst_7_1_N0 ), .Z(n1871) );
  OR2 U2021 ( .A(n1873), .B(AddKeyConstXOR_XORInst_7_3_N0 ), .Z(n1869) );
  BIC2 U2022 ( .A(n1852), .B(AddKeyConstXOR_XORInst_7_1_N0 ), .Z(n1873) );
  ORN2 U2023 ( .A(n1874), .B(AddKeyConstXOR_XORInst_7_2_N0 ), .Z(n1852) );
  ORN2 U2024 ( .A(n1678), .B(n1273), .Z(n1866) );
  BIC2 U2025 ( .A(n1875), .B(n1876), .Z(n1678) );
  AND2 U2026 ( .A(n1877), .B(n1830), .Z(n1876) );
  NOT1 U2027 ( .A(AddKeyConstXOR_XORInst_3_2_N0 ), .Z(n1830) );
  OR2 U2028 ( .A(n1841), .B(AddKeyConstXOR_XORInst_3_1_N0 ), .Z(n1877) );
  AND2 U2029 ( .A(AddKeyConstXOR_XORInst_3_3_N0 ), .B(
        AddKeyConstXOR_XORInst_3_0_N1 ), .Z(n1841) );
  OR2 U2030 ( .A(n1878), .B(AddKeyConstXOR_XORInst_3_3_N0 ), .Z(n1875) );
  BIC2 U2031 ( .A(n1861), .B(AddKeyConstXOR_XORInst_3_1_N0 ), .Z(n1878) );
  ORN2 U2032 ( .A(n1831), .B(AddKeyConstXOR_XORInst_3_2_N0 ), .Z(n1861) );
  AND2 U2033 ( .A(Plaintext[12]), .B(rst), .Z(n1864) );
  ORN2 U2034 ( .A(n1879), .B(n1880), .Z(StateRegInput[11]) );
  AND2 U2035 ( .A(n1881), .B(n1882), .Z(n1880) );
  ORN2 U2036 ( .A(n1249), .B(n1883), .Z(n1882) );
  XOR2 U2037 ( .A(n1826), .B(n1511), .Z(n1883) );
  BIC2 U2038 ( .A(n1884), .B(n1885), .Z(n1511) );
  BIC2 U2039 ( .A(n1886), .B(AddKeyConstXOR_XORInst_8_3_N0 ), .Z(n1885) );
  ORN2 U2040 ( .A(n1746), .B(AddKeyConstXOR_XORInst_8_1_N0 ), .Z(n1886) );
  ORN2 U2041 ( .A(AddKeyConstXOR_XORInst_8_2_N0 ), .B(n1887), .Z(n1884) );
  NOT1 U2042 ( .A(AddKeyConstXOR_XORInst_8_1_N0 ), .Z(n1887) );
  XOR2 U2043 ( .A(n1360), .B(n1271), .Z(n1826) );
  BIC2 U2044 ( .A(n1888), .B(n1889), .Z(n1271) );
  AND2 U2045 ( .A(AddKeyConstXOR_XORInst_7_1_N0 ), .B(n1890), .Z(n1889) );
  ORN2 U2046 ( .A(n1855), .B(AddKeyConstXOR_XORInst_7_3_N0 ), .Z(n1888) );
  ORN2 U2047 ( .A(n1891), .B(n1892), .Z(n1360) );
  ORN2 U2048 ( .A(n1858), .B(AddKeyConstXOR_XORInst_13_3_N0 ), .Z(n1892) );
  AND2 U2049 ( .A(AddKeyConstXOR_XORInst_13_1_N0 ), .B(n1893), .Z(n1891) );
  ORN2 U2050 ( .A(n1254), .B(n1512), .Z(n1881) );
  BIC2 U2051 ( .A(n1894), .B(n1895), .Z(n1512) );
  AND2 U2052 ( .A(AddKeyConstXOR_XORInst_2_1_N0 ), .B(n1896), .Z(n1895) );
  ORN2 U2053 ( .A(n1851), .B(AddKeyConstXOR_XORInst_2_3_N0 ), .Z(n1894) );
  AND2 U2054 ( .A(Plaintext[11]), .B(rst), .Z(n1879) );
  ORN2 U2055 ( .A(n1897), .B(n1898), .Z(StateRegInput[10]) );
  AND2 U2056 ( .A(n1899), .B(n1900), .Z(n1898) );
  ORN2 U2057 ( .A(n1249), .B(n1901), .Z(n1900) );
  XOR2 U2058 ( .A(n1837), .B(n1590), .Z(n1901) );
  BIC2 U2059 ( .A(n1902), .B(n1903), .Z(n1590) );
  AND2 U2060 ( .A(n1904), .B(AddKeyConstXOR_XORInst_8_1_N0 ), .Z(n1903) );
  ORN2 U2061 ( .A(n1905), .B(n1744), .Z(n1904) );
  NOT1 U2062 ( .A(AddKeyConstXOR_XORInst_8_2_N0 ), .Z(n1744) );
  AND2 U2063 ( .A(AddKeyConstXOR_XORInst_8_3_N0 ), .B(
        AddKeyConstXOR_XORInst_8_0_N1 ), .Z(n1905) );
  OR2 U2064 ( .A(AddKeyConstXOR_XORInst_8_3_N0 ), .B(
        AddKeyConstXOR_XORInst_8_0_N1 ), .Z(n1902) );
  XOR2 U2065 ( .A(n1367), .B(n1280), .Z(n1837) );
  BIC2 U2066 ( .A(n1890), .B(n1906), .Z(n1280) );
  AND2 U2067 ( .A(AddKeyConstXOR_XORInst_7_1_N0 ), .B(n1907), .Z(n1906) );
  ORN2 U2068 ( .A(n1872), .B(n1855), .Z(n1907) );
  NOT1 U2069 ( .A(AddKeyConstXOR_XORInst_7_2_N0 ), .Z(n1855) );
  AND2 U2070 ( .A(AddKeyConstXOR_XORInst_7_3_N0 ), .B(
        AddKeyConstXOR_XORInst_7_0_N1 ), .Z(n1872) );
  OR2 U2071 ( .A(AddKeyConstXOR_XORInst_7_3_N0 ), .B(
        AddKeyConstXOR_XORInst_7_0_N1 ), .Z(n1890) );
  ORN2 U2072 ( .A(n1908), .B(n1893), .Z(n1367) );
  ORN2 U2073 ( .A(AddKeyConstXOR_XORInst_13_0_N1 ), .B(n1909), .Z(n1893) );
  AND2 U2074 ( .A(AddKeyConstXOR_XORInst_13_1_N0 ), .B(n1910), .Z(n1908) );
  ORN2 U2075 ( .A(n1911), .B(n1858), .Z(n1910) );
  AND2 U2076 ( .A(AddKeyConstXOR_XORInst_13_3_N0 ), .B(
        AddKeyConstXOR_XORInst_13_0_N1 ), .Z(n1911) );
  ORN2 U2077 ( .A(n1634), .B(n1273), .Z(n1899) );
  BIC2 U2078 ( .A(n1896), .B(n1912), .Z(n1634) );
  AND2 U2079 ( .A(AddKeyConstXOR_XORInst_2_1_N0 ), .B(n1913), .Z(n1912) );
  ORN2 U2080 ( .A(n1914), .B(n1851), .Z(n1913) );
  AND2 U2081 ( .A(AddKeyConstXOR_XORInst_2_3_N0 ), .B(
        AddKeyConstXOR_XORInst_2_0_N1 ), .Z(n1914) );
  ORN2 U2082 ( .A(AddKeyConstXOR_XORInst_2_0_N1 ), .B(n1915), .Z(n1896) );
  AND2 U2083 ( .A(Plaintext[10]), .B(rst), .Z(n1897) );
  ORN2 U2084 ( .A(n1916), .B(n1917), .Z(StateRegInput[0]) );
  AND2 U2085 ( .A(n1918), .B(n1919), .Z(n1917) );
  ORN2 U2086 ( .A(n1249), .B(n1920), .Z(n1919) );
  XOR2 U2087 ( .A(n1407), .B(n1381), .Z(n1920) );
  BIC2 U2088 ( .A(n1921), .B(n1922), .Z(n1381) );
  AND2 U2089 ( .A(n1923), .B(AddKeyConstXOR_XORInst_13_0_N1 ), .Z(n1922) );
  XOR2 U2090 ( .A(n1858), .B(n1909), .Z(n1923) );
  NOT1 U2091 ( .A(AddKeyConstXOR_XORInst_13_3_N0 ), .Z(n1909) );
  NOT1 U2092 ( .A(AddKeyConstXOR_XORInst_13_2_N0 ), .Z(n1858) );
  ORN2 U2093 ( .A(n1924), .B(AddKeyConstXOR_XORInst_13_1_N0 ), .Z(n1921) );
  AND2 U2094 ( .A(AddKeyConstXOR_XORInst_13_3_N0 ), .B(
        AddKeyConstXOR_XORInst_13_2_N0 ), .Z(n1924) );
  XOR2 U2095 ( .A(n1264), .B(n1263), .Z(n1407) );
  BIC2 U2096 ( .A(n1925), .B(n1926), .Z(n1263) );
  AND2 U2097 ( .A(n1927), .B(AddKeyConstXOR_XORInst_8_0_N1 ), .Z(n1926) );
  XOR2 U2098 ( .A(AddKeyConstXOR_XORInst_8_2_N0 ), .B(
        AddKeyConstXOR_XORInst_8_3_N0 ), .Z(n1927) );
  ORN2 U2099 ( .A(n1928), .B(AddKeyConstXOR_XORInst_8_1_N0 ), .Z(n1925) );
  AND2 U2100 ( .A(AddKeyConstXOR_XORInst_8_3_N0 ), .B(
        AddKeyConstXOR_XORInst_8_2_N0 ), .Z(n1928) );
  ORN2 U2101 ( .A(n1929), .B(n1930), .Z(n1264) );
  ORN2 U2102 ( .A(n1931), .B(AddKeyConstXOR_XORInst_2_1_N0 ), .Z(n1930) );
  AND2 U2103 ( .A(AddKeyConstXOR_XORInst_2_3_N0 ), .B(
        AddKeyConstXOR_XORInst_2_2_N0 ), .Z(n1931) );
  AND2 U2104 ( .A(n1932), .B(AddKeyConstXOR_XORInst_2_0_N1 ), .Z(n1929) );
  XOR2 U2105 ( .A(n1851), .B(n1915), .Z(n1932) );
  NOT1 U2106 ( .A(AddKeyConstXOR_XORInst_2_3_N0 ), .Z(n1915) );
  NOT1 U2107 ( .A(AddKeyConstXOR_XORInst_2_2_N0 ), .Z(n1851) );
  OR2 U2108 ( .A(rst), .B(n1933), .Z(n1249) );
  ORN2 U2109 ( .A(n1351), .B(n1273), .Z(n1918) );
  BIC2 U2110 ( .A(n1934), .B(n1935), .Z(n1351) );
  AND2 U2111 ( .A(n1936), .B(n1516), .Z(n1935) );
  NOT1 U2112 ( .A(AddKeyConstXOR_XORInst_0_2_N0 ), .Z(n1516) );
  OR2 U2113 ( .A(n1638), .B(AddKeyConstXOR_XORInst_0_1_N0 ), .Z(n1936) );
  AND2 U2114 ( .A(AddKeyConstXOR_XORInst_0_3_N0 ), .B(
        AddKeyConstXOR_XORInst_0_0_N1 ), .Z(n1638) );
  OR2 U2115 ( .A(n1937), .B(AddKeyConstXOR_XORInst_0_3_N0 ), .Z(n1934) );
  BIC2 U2116 ( .A(n1747), .B(AddKeyConstXOR_XORInst_0_1_N0 ), .Z(n1937) );
  ORN2 U2117 ( .A(n1517), .B(AddKeyConstXOR_XORInst_0_2_N0 ), .Z(n1747) );
  AND2 U2118 ( .A(Plaintext[0]), .B(rst), .Z(n1916) );
  ORN2 U2119 ( .A(n1938), .B(n1254), .Z(FSMSelected[4]) );
  NOT1 U2120 ( .A(n1273), .Z(n1254) );
  AND2 U2121 ( .A(n1933), .B(n1939), .Z(n1273) );
  BIC2 U2122 ( .A(FSM[4] ), .B(rst), .Z(n1938) );
  AND2 U2123 ( .A(n1940), .B(n1939), .Z(FSMSelected[3]) );
  ORN2 U2124 ( .A(n1941), .B(n1942), .Z(n1940) );
  ORN2 U2125 ( .A(n1943), .B(n1944), .Z(n1942) );
  BIC2 U2126 ( .A(Round[3]), .B(n1945), .Z(n1941) );
  AND2 U2127 ( .A(n1944), .B(n1946), .Z(n1945) );
  AND2 U2128 ( .A(n1947), .B(n1939), .Z(FSMSelected[2]) );
  ORN2 U2129 ( .A(n1948), .B(n1949), .Z(n1947) );
  AND2 U2130 ( .A(n1950), .B(n1951), .Z(n1949) );
  ORN2 U2131 ( .A(n1944), .B(n1946), .Z(n1951) );
  AND2 U2132 ( .A(Round[1]), .B(n1952), .Z(n1944) );
  ORN2 U2133 ( .A(FSM[4] ), .B(n1953), .Z(n1950) );
  ORN2 U2134 ( .A(n1954), .B(n1955), .Z(n1948) );
  AND2 U2135 ( .A(n1956), .B(n1939), .Z(FSMSelected[1]) );
  ORN2 U2136 ( .A(n1957), .B(n1958), .Z(n1956) );
  AND2 U2137 ( .A(n1959), .B(n1960), .Z(n1958) );
  ORN2 U2138 ( .A(n1961), .B(n1962), .Z(n1957) );
  ORN2 U2139 ( .A(n1952), .B(Round[1]), .Z(n1962) );
  NOT1 U2140 ( .A(FSM[4] ), .Z(n1952) );
  AND2 U2141 ( .A(n1963), .B(n1964), .Z(n1961) );
  BIC2 U2142 ( .A(Round[0]), .B(FSM[4] ), .Z(n1963) );
  AND2 U2143 ( .A(n1965), .B(n1939), .Z(FSMSelected[0]) );
  NOT1 U2144 ( .A(rst), .Z(n1939) );
  ORN2 U2145 ( .A(n1966), .B(n1967), .Z(n1965) );
  AND2 U2146 ( .A(n1968), .B(n1955), .Z(n1967) );
  ORN2 U2147 ( .A(FSM[4] ), .B(n1959), .Z(n1966) );
  XOR2 U2148 ( .A(n1969), .B(StateRegOutput[39]), .Z(
        AddKeyConstXOR_XORInst_9_3_N0 ) );
  ORN2 U2149 ( .A(n1970), .B(n1971), .Z(n1969) );
  ORN2 U2150 ( .A(n1972), .B(Key[39]), .Z(n1971) );
  BIC2 U2151 ( .A(n1973), .B(n1974), .Z(n1972) );
  OR2 U2152 ( .A(Key[103]), .B(n1975), .Z(n1973) );
  AND2 U2153 ( .A(n1976), .B(Key[103]), .Z(n1970) );
  ORN2 U2154 ( .A(n1977), .B(n1978), .Z(n1976) );
  BIC2 U2155 ( .A(n1979), .B(Key[39]), .Z(n1977) );
  XOR2 U2156 ( .A(n1980), .B(StateRegOutput[38]), .Z(
        AddKeyConstXOR_XORInst_9_2_N0 ) );
  ORN2 U2157 ( .A(n1981), .B(n1982), .Z(n1980) );
  ORN2 U2158 ( .A(n1983), .B(Key[38]), .Z(n1982) );
  BIC2 U2159 ( .A(n1984), .B(n1974), .Z(n1983) );
  OR2 U2160 ( .A(Key[102]), .B(n1975), .Z(n1984) );
  AND2 U2161 ( .A(n1985), .B(Key[102]), .Z(n1981) );
  ORN2 U2162 ( .A(n1986), .B(n1978), .Z(n1985) );
  BIC2 U2163 ( .A(n1979), .B(Key[38]), .Z(n1986) );
  XOR2 U2164 ( .A(n1987), .B(StateRegOutput[37]), .Z(
        AddKeyConstXOR_XORInst_9_1_N0 ) );
  ORN2 U2165 ( .A(n1988), .B(n1989), .Z(n1987) );
  ORN2 U2166 ( .A(n1990), .B(Key[37]), .Z(n1989) );
  BIC2 U2167 ( .A(n1991), .B(n1974), .Z(n1990) );
  OR2 U2168 ( .A(Key[101]), .B(n1975), .Z(n1991) );
  AND2 U2169 ( .A(n1992), .B(Key[101]), .Z(n1988) );
  ORN2 U2170 ( .A(n1993), .B(n1978), .Z(n1992) );
  BIC2 U2171 ( .A(n1979), .B(Key[37]), .Z(n1993) );
  NOT1 U2172 ( .A(n1698), .Z(AddKeyConstXOR_XORInst_9_0_N1 ) );
  XOR2 U2173 ( .A(n1994), .B(n1995), .Z(n1698) );
  AND2 U2174 ( .A(n1996), .B(n1997), .Z(n1995) );
  ORN2 U2175 ( .A(n1964), .B(n1946), .Z(n1997) );
  AND2 U2176 ( .A(n1955), .B(n1998), .Z(n1996) );
  XOR2 U2177 ( .A(n1999), .B(StateRegOutput[36]), .Z(n1994) );
  ORN2 U2178 ( .A(n2000), .B(n2001), .Z(n1999) );
  ORN2 U2179 ( .A(n2002), .B(n2003), .Z(n2001) );
  AND2 U2180 ( .A(n2004), .B(n2005), .Z(n2003) );
  ORN2 U2181 ( .A(n1974), .B(Key[100]), .Z(n2004) );
  AND2 U2182 ( .A(Key[100]), .B(n2006), .Z(n2000) );
  ORN2 U2183 ( .A(n2007), .B(n1978), .Z(n2006) );
  BIC2 U2184 ( .A(n2002), .B(n1975), .Z(n2007) );
  NOT1 U2185 ( .A(Key[36]), .Z(n2002) );
  XOR2 U2186 ( .A(n2008), .B(StateRegOutput[35]), .Z(
        AddKeyConstXOR_XORInst_8_3_N0 ) );
  ORN2 U2187 ( .A(n2009), .B(n2010), .Z(n2008) );
  ORN2 U2188 ( .A(n2011), .B(Key[99]), .Z(n2010) );
  AND2 U2189 ( .A(n2012), .B(n1978), .Z(n2011) );
  OR2 U2190 ( .A(Key[35]), .B(n1975), .Z(n2012) );
  AND2 U2191 ( .A(n2013), .B(Key[35]), .Z(n2009) );
  OR2 U2192 ( .A(n2014), .B(n1974), .Z(n2013) );
  BIC2 U2193 ( .A(n1979), .B(Key[99]), .Z(n2014) );
  XOR2 U2194 ( .A(n2015), .B(StateRegOutput[34]), .Z(
        AddKeyConstXOR_XORInst_8_2_N0 ) );
  ORN2 U2195 ( .A(n2016), .B(n2017), .Z(n2015) );
  ORN2 U2196 ( .A(n2018), .B(Key[98]), .Z(n2017) );
  AND2 U2197 ( .A(n2019), .B(n1978), .Z(n2018) );
  OR2 U2198 ( .A(Key[34]), .B(n1975), .Z(n2019) );
  AND2 U2199 ( .A(n2020), .B(Key[34]), .Z(n2016) );
  OR2 U2200 ( .A(n2021), .B(n1974), .Z(n2020) );
  BIC2 U2201 ( .A(n1979), .B(Key[98]), .Z(n2021) );
  XOR2 U2202 ( .A(n2022), .B(StateRegOutput[33]), .Z(
        AddKeyConstXOR_XORInst_8_1_N0 ) );
  ORN2 U2203 ( .A(n2023), .B(n2024), .Z(n2022) );
  ORN2 U2204 ( .A(n2025), .B(Key[97]), .Z(n2024) );
  AND2 U2205 ( .A(n2026), .B(n1978), .Z(n2025) );
  OR2 U2206 ( .A(Key[33]), .B(n1975), .Z(n2026) );
  AND2 U2207 ( .A(n2027), .B(Key[33]), .Z(n2023) );
  OR2 U2208 ( .A(n2028), .B(n1974), .Z(n2027) );
  BIC2 U2209 ( .A(n1979), .B(Key[97]), .Z(n2028) );
  NOT1 U2210 ( .A(n1746), .Z(AddKeyConstXOR_XORInst_8_0_N1 ) );
  XOR2 U2211 ( .A(n2029), .B(n2030), .Z(n1746) );
  AND2 U2212 ( .A(n2031), .B(n2032), .Z(n2030) );
  AND2 U2213 ( .A(n2033), .B(n2034), .Z(n2032) );
  ORN2 U2214 ( .A(n2035), .B(n2036), .Z(n2033) );
  AND2 U2215 ( .A(n2037), .B(n1959), .Z(n2035) );
  AND2 U2216 ( .A(n2038), .B(n2039), .Z(n2031) );
  ORN2 U2217 ( .A(n1978), .B(n2040), .Z(n2038) );
  XOR2 U2218 ( .A(n2041), .B(StateRegOutput[32]), .Z(n2029) );
  ORN2 U2219 ( .A(n2042), .B(n2043), .Z(n2041) );
  ORN2 U2220 ( .A(n2044), .B(n2045), .Z(n2043) );
  BIC2 U2221 ( .A(n2046), .B(n1974), .Z(n2045) );
  ORN2 U2222 ( .A(Round[0]), .B(Key[32]), .Z(n2046) );
  AND2 U2223 ( .A(Key[32]), .B(n2047), .Z(n2042) );
  OR2 U2224 ( .A(n2048), .B(n1974), .Z(n2047) );
  BIC2 U2225 ( .A(n2044), .B(n1975), .Z(n2048) );
  NOT1 U2226 ( .A(Key[96]), .Z(n2044) );
  XOR2 U2227 ( .A(n2049), .B(StateRegOutput[31]), .Z(
        AddKeyConstXOR_XORInst_7_3_N0 ) );
  ORN2 U2228 ( .A(n2050), .B(n2051), .Z(n2049) );
  ORN2 U2229 ( .A(n2052), .B(Key[95]), .Z(n2051) );
  AND2 U2230 ( .A(n2053), .B(n1978), .Z(n2052) );
  OR2 U2231 ( .A(Key[31]), .B(n1975), .Z(n2053) );
  AND2 U2232 ( .A(n2054), .B(Key[31]), .Z(n2050) );
  OR2 U2233 ( .A(n2055), .B(n1974), .Z(n2054) );
  BIC2 U2234 ( .A(n1979), .B(Key[95]), .Z(n2055) );
  XOR2 U2235 ( .A(n2056), .B(StateRegOutput[30]), .Z(
        AddKeyConstXOR_XORInst_7_2_N0 ) );
  ORN2 U2236 ( .A(n2057), .B(n2058), .Z(n2056) );
  ORN2 U2237 ( .A(n2059), .B(Key[94]), .Z(n2058) );
  AND2 U2238 ( .A(n2060), .B(n1978), .Z(n2059) );
  OR2 U2239 ( .A(Key[30]), .B(n1975), .Z(n2060) );
  AND2 U2240 ( .A(n2061), .B(Key[30]), .Z(n2057) );
  OR2 U2241 ( .A(n2062), .B(n1974), .Z(n2061) );
  BIC2 U2242 ( .A(n1979), .B(Key[94]), .Z(n2062) );
  XOR2 U2243 ( .A(n2063), .B(StateRegOutput[29]), .Z(
        AddKeyConstXOR_XORInst_7_1_N0 ) );
  ORN2 U2244 ( .A(n2064), .B(n2065), .Z(n2063) );
  ORN2 U2245 ( .A(n2066), .B(Key[93]), .Z(n2065) );
  AND2 U2246 ( .A(n2067), .B(n1978), .Z(n2066) );
  OR2 U2247 ( .A(Key[29]), .B(n1975), .Z(n2067) );
  AND2 U2248 ( .A(n2068), .B(Key[29]), .Z(n2064) );
  OR2 U2249 ( .A(n2069), .B(n1974), .Z(n2068) );
  BIC2 U2250 ( .A(n1979), .B(Key[93]), .Z(n2069) );
  NOT1 U2251 ( .A(n1874), .Z(AddKeyConstXOR_XORInst_7_0_N1 ) );
  XOR2 U2252 ( .A(n2070), .B(n2071), .Z(n1874) );
  AND2 U2253 ( .A(n2072), .B(n2073), .Z(n2071) );
  AND2 U2254 ( .A(n2037), .B(n2074), .Z(n2073) );
  AND2 U2255 ( .A(n2075), .B(n1960), .Z(n2072) );
  XOR2 U2256 ( .A(n2076), .B(StateRegOutput[28]), .Z(n2070) );
  ORN2 U2257 ( .A(n2077), .B(n2078), .Z(n2076) );
  ORN2 U2258 ( .A(n2079), .B(n2080), .Z(n2078) );
  BIC2 U2259 ( .A(n2081), .B(n1974), .Z(n2080) );
  ORN2 U2260 ( .A(Round[0]), .B(Key[28]), .Z(n2081) );
  AND2 U2261 ( .A(Key[28]), .B(n2082), .Z(n2077) );
  OR2 U2262 ( .A(n2083), .B(n1974), .Z(n2082) );
  BIC2 U2263 ( .A(n2079), .B(n1975), .Z(n2083) );
  NOT1 U2264 ( .A(Key[92]), .Z(n2079) );
  XOR2 U2265 ( .A(n2084), .B(StateRegOutput[27]), .Z(
        AddKeyConstXOR_XORInst_6_3_N0 ) );
  ORN2 U2266 ( .A(n2085), .B(n2086), .Z(n2084) );
  ORN2 U2267 ( .A(n2087), .B(Key[91]), .Z(n2086) );
  AND2 U2268 ( .A(n2088), .B(n1978), .Z(n2087) );
  OR2 U2269 ( .A(Key[27]), .B(n1975), .Z(n2088) );
  AND2 U2270 ( .A(n2089), .B(Key[27]), .Z(n2085) );
  OR2 U2271 ( .A(n2090), .B(n1974), .Z(n2089) );
  BIC2 U2272 ( .A(n1979), .B(Key[91]), .Z(n2090) );
  XOR2 U2273 ( .A(n2091), .B(StateRegOutput[26]), .Z(
        AddKeyConstXOR_XORInst_6_2_N0 ) );
  ORN2 U2274 ( .A(n2092), .B(n2093), .Z(n2091) );
  ORN2 U2275 ( .A(n2094), .B(Key[90]), .Z(n2093) );
  AND2 U2276 ( .A(n2095), .B(n1978), .Z(n2094) );
  OR2 U2277 ( .A(Key[26]), .B(n1975), .Z(n2095) );
  AND2 U2278 ( .A(n2096), .B(Key[26]), .Z(n2092) );
  OR2 U2279 ( .A(n2097), .B(n1974), .Z(n2096) );
  BIC2 U2280 ( .A(n1979), .B(Key[90]), .Z(n2097) );
  XOR2 U2281 ( .A(n2098), .B(StateRegOutput[25]), .Z(
        AddKeyConstXOR_XORInst_6_1_N0 ) );
  ORN2 U2282 ( .A(n2099), .B(n2100), .Z(n2098) );
  ORN2 U2283 ( .A(n2101), .B(Key[89]), .Z(n2100) );
  AND2 U2284 ( .A(n2102), .B(n1978), .Z(n2101) );
  OR2 U2285 ( .A(Key[25]), .B(n1975), .Z(n2102) );
  AND2 U2286 ( .A(n2103), .B(Key[25]), .Z(n2099) );
  OR2 U2287 ( .A(n2104), .B(n1974), .Z(n2103) );
  BIC2 U2288 ( .A(n1979), .B(Key[89]), .Z(n2104) );
  NOT1 U2289 ( .A(n1770), .Z(AddKeyConstXOR_XORInst_6_0_N1 ) );
  XOR2 U2290 ( .A(n2105), .B(n2106), .Z(n1770) );
  AND2 U2291 ( .A(n2107), .B(n2108), .Z(n2106) );
  AND2 U2292 ( .A(n2034), .B(n1943), .Z(n2107) );
  XOR2 U2293 ( .A(n2109), .B(StateRegOutput[24]), .Z(n2105) );
  ORN2 U2294 ( .A(n2110), .B(n2111), .Z(n2109) );
  ORN2 U2295 ( .A(n2112), .B(n2113), .Z(n2111) );
  BIC2 U2296 ( .A(n2114), .B(n1974), .Z(n2113) );
  ORN2 U2297 ( .A(Round[0]), .B(Key[24]), .Z(n2114) );
  AND2 U2298 ( .A(Key[24]), .B(n2115), .Z(n2110) );
  OR2 U2299 ( .A(n2116), .B(n1974), .Z(n2115) );
  BIC2 U2300 ( .A(n2112), .B(n1975), .Z(n2116) );
  NOT1 U2301 ( .A(Key[88]), .Z(n2112) );
  XOR2 U2302 ( .A(n2117), .B(StateRegOutput[23]), .Z(
        AddKeyConstXOR_XORInst_5_3_N0 ) );
  ORN2 U2303 ( .A(n2118), .B(n2119), .Z(n2117) );
  ORN2 U2304 ( .A(n2120), .B(Key[87]), .Z(n2119) );
  AND2 U2305 ( .A(n2121), .B(n1978), .Z(n2120) );
  OR2 U2306 ( .A(Key[23]), .B(n1975), .Z(n2121) );
  AND2 U2307 ( .A(n2122), .B(Key[23]), .Z(n2118) );
  OR2 U2308 ( .A(n2123), .B(n1974), .Z(n2122) );
  BIC2 U2309 ( .A(n1979), .B(Key[87]), .Z(n2123) );
  XOR2 U2310 ( .A(n2124), .B(StateRegOutput[22]), .Z(
        AddKeyConstXOR_XORInst_5_2_N0 ) );
  ORN2 U2311 ( .A(n2125), .B(n2126), .Z(n2124) );
  ORN2 U2312 ( .A(n2127), .B(Key[86]), .Z(n2126) );
  AND2 U2313 ( .A(n2128), .B(n1978), .Z(n2127) );
  OR2 U2314 ( .A(Key[22]), .B(n1975), .Z(n2128) );
  AND2 U2315 ( .A(n2129), .B(Key[22]), .Z(n2125) );
  OR2 U2316 ( .A(n2130), .B(n1974), .Z(n2129) );
  BIC2 U2317 ( .A(n1979), .B(Key[86]), .Z(n2130) );
  XOR2 U2318 ( .A(n2131), .B(StateRegOutput[21]), .Z(
        AddKeyConstXOR_XORInst_5_1_N0 ) );
  ORN2 U2319 ( .A(n2132), .B(n2133), .Z(n2131) );
  ORN2 U2320 ( .A(n2134), .B(Key[85]), .Z(n2133) );
  AND2 U2321 ( .A(n2135), .B(n1978), .Z(n2134) );
  OR2 U2322 ( .A(Key[21]), .B(n1975), .Z(n2135) );
  AND2 U2323 ( .A(n2136), .B(Key[21]), .Z(n2132) );
  OR2 U2324 ( .A(n2137), .B(n1974), .Z(n2136) );
  BIC2 U2325 ( .A(n1979), .B(Key[85]), .Z(n2137) );
  NOT1 U2326 ( .A(n1703), .Z(AddKeyConstXOR_XORInst_5_0_N1 ) );
  XOR2 U2327 ( .A(n2138), .B(n2139), .Z(n1703) );
  AND2 U2328 ( .A(n2140), .B(n2141), .Z(n2139) );
  BIC2 U2329 ( .A(n2142), .B(n2143), .Z(n2141) );
  ORN2 U2330 ( .A(n2144), .B(n2145), .Z(n2142) );
  AND2 U2331 ( .A(n2146), .B(n2147), .Z(n2140) );
  ORN2 U2332 ( .A(n2036), .B(n2148), .Z(n2147) );
  ORN2 U2333 ( .A(Round[1]), .B(n2149), .Z(n2146) );
  XOR2 U2334 ( .A(n2150), .B(StateRegOutput[20]), .Z(n2138) );
  ORN2 U2335 ( .A(n2151), .B(n2152), .Z(n2150) );
  ORN2 U2336 ( .A(n2153), .B(n2154), .Z(n2152) );
  BIC2 U2337 ( .A(n2155), .B(n1974), .Z(n2154) );
  ORN2 U2338 ( .A(Round[0]), .B(Key[20]), .Z(n2155) );
  AND2 U2339 ( .A(Key[20]), .B(n2156), .Z(n2151) );
  OR2 U2340 ( .A(n2157), .B(n1974), .Z(n2156) );
  BIC2 U2341 ( .A(n2153), .B(n1975), .Z(n2157) );
  NOT1 U2342 ( .A(Key[84]), .Z(n2153) );
  XOR2 U2343 ( .A(n2158), .B(StateRegOutput[19]), .Z(
        AddKeyConstXOR_XORInst_4_3_N0 ) );
  ORN2 U2344 ( .A(n2159), .B(n2160), .Z(n2158) );
  ORN2 U2345 ( .A(n2161), .B(Key[83]), .Z(n2160) );
  AND2 U2346 ( .A(n2162), .B(n1978), .Z(n2161) );
  OR2 U2347 ( .A(Key[19]), .B(n1975), .Z(n2162) );
  AND2 U2348 ( .A(n2163), .B(Key[19]), .Z(n2159) );
  OR2 U2349 ( .A(n2164), .B(n1974), .Z(n2163) );
  BIC2 U2350 ( .A(n1979), .B(Key[83]), .Z(n2164) );
  XOR2 U2351 ( .A(n2165), .B(StateRegOutput[18]), .Z(
        AddKeyConstXOR_XORInst_4_2_N0 ) );
  ORN2 U2352 ( .A(n2166), .B(n2167), .Z(n2165) );
  ORN2 U2353 ( .A(n2168), .B(Key[82]), .Z(n2167) );
  AND2 U2354 ( .A(n2169), .B(n1978), .Z(n2168) );
  OR2 U2355 ( .A(Key[18]), .B(n1975), .Z(n2169) );
  AND2 U2356 ( .A(n2170), .B(Key[18]), .Z(n2166) );
  OR2 U2357 ( .A(n2171), .B(n1974), .Z(n2170) );
  BIC2 U2358 ( .A(n1979), .B(Key[82]), .Z(n2171) );
  XOR2 U2359 ( .A(n2172), .B(StateRegOutput[17]), .Z(
        AddKeyConstXOR_XORInst_4_1_N0 ) );
  ORN2 U2360 ( .A(n2173), .B(n2174), .Z(n2172) );
  ORN2 U2361 ( .A(n2175), .B(Key[81]), .Z(n2174) );
  AND2 U2362 ( .A(n2176), .B(n1978), .Z(n2175) );
  OR2 U2363 ( .A(Key[17]), .B(n1975), .Z(n2176) );
  AND2 U2364 ( .A(n2177), .B(Key[17]), .Z(n2173) );
  OR2 U2365 ( .A(n2178), .B(n1974), .Z(n2177) );
  BIC2 U2366 ( .A(n1979), .B(Key[81]), .Z(n2178) );
  NOT1 U2367 ( .A(n1780), .Z(AddKeyConstXOR_XORInst_4_0_N1 ) );
  XOR2 U2368 ( .A(n2179), .B(n2180), .Z(n1780) );
  AND2 U2369 ( .A(n2181), .B(n2182), .Z(n2180) );
  BIC2 U2370 ( .A(n2183), .B(n2143), .Z(n2182) );
  AND2 U2371 ( .A(n2184), .B(n2039), .Z(n2181) );
  ORN2 U2372 ( .A(Round[2]), .B(n2040), .Z(n2184) );
  XOR2 U2373 ( .A(n2185), .B(StateRegOutput[16]), .Z(n2179) );
  ORN2 U2374 ( .A(n2186), .B(n2187), .Z(n2185) );
  ORN2 U2375 ( .A(n2188), .B(n2189), .Z(n2187) );
  BIC2 U2376 ( .A(n2190), .B(n1974), .Z(n2189) );
  ORN2 U2377 ( .A(Round[0]), .B(Key[16]), .Z(n2190) );
  AND2 U2378 ( .A(Key[16]), .B(n2191), .Z(n2186) );
  OR2 U2379 ( .A(n2192), .B(n1974), .Z(n2191) );
  BIC2 U2380 ( .A(n2188), .B(n1975), .Z(n2192) );
  NOT1 U2381 ( .A(Key[80]), .Z(n2188) );
  XOR2 U2382 ( .A(n2193), .B(StateRegOutput[15]), .Z(
        AddKeyConstXOR_XORInst_3_3_N0 ) );
  ORN2 U2383 ( .A(n2194), .B(n2195), .Z(n2193) );
  ORN2 U2384 ( .A(n2196), .B(Key[79]), .Z(n2195) );
  AND2 U2385 ( .A(n2197), .B(n1978), .Z(n2196) );
  OR2 U2386 ( .A(Key[15]), .B(n1975), .Z(n2197) );
  AND2 U2387 ( .A(n2198), .B(Key[15]), .Z(n2194) );
  OR2 U2388 ( .A(n2199), .B(n1974), .Z(n2198) );
  BIC2 U2389 ( .A(n1979), .B(Key[79]), .Z(n2199) );
  XOR2 U2390 ( .A(n2200), .B(StateRegOutput[14]), .Z(
        AddKeyConstXOR_XORInst_3_2_N0 ) );
  ORN2 U2391 ( .A(n2201), .B(n2202), .Z(n2200) );
  ORN2 U2392 ( .A(n2203), .B(Key[78]), .Z(n2202) );
  AND2 U2393 ( .A(n2204), .B(n1978), .Z(n2203) );
  OR2 U2394 ( .A(Key[14]), .B(n1975), .Z(n2204) );
  AND2 U2395 ( .A(n2205), .B(Key[14]), .Z(n2201) );
  OR2 U2396 ( .A(n2206), .B(n1974), .Z(n2205) );
  BIC2 U2397 ( .A(n1979), .B(Key[78]), .Z(n2206) );
  XOR2 U2398 ( .A(n2207), .B(StateRegOutput[13]), .Z(
        AddKeyConstXOR_XORInst_3_1_N0 ) );
  ORN2 U2399 ( .A(n2208), .B(n2209), .Z(n2207) );
  ORN2 U2400 ( .A(n2210), .B(Key[77]), .Z(n2209) );
  AND2 U2401 ( .A(n2211), .B(n1978), .Z(n2210) );
  OR2 U2402 ( .A(Key[13]), .B(n1975), .Z(n2211) );
  AND2 U2403 ( .A(n2212), .B(Key[13]), .Z(n2208) );
  OR2 U2404 ( .A(n2213), .B(n1974), .Z(n2212) );
  BIC2 U2405 ( .A(n1979), .B(Key[77]), .Z(n2213) );
  NOT1 U2406 ( .A(n1831), .Z(AddKeyConstXOR_XORInst_3_0_N1 ) );
  XOR2 U2407 ( .A(n2214), .B(n2215), .Z(n1831) );
  AND2 U2408 ( .A(n2216), .B(n2075), .Z(n2215) );
  ORN2 U2409 ( .A(Round[1]), .B(n2217), .Z(n2216) );
  XOR2 U2410 ( .A(n2218), .B(StateRegOutput[12]), .Z(n2214) );
  ORN2 U2411 ( .A(n2219), .B(n2220), .Z(n2218) );
  ORN2 U2412 ( .A(n2221), .B(n2222), .Z(n2220) );
  BIC2 U2413 ( .A(n2223), .B(n1974), .Z(n2222) );
  ORN2 U2414 ( .A(Round[0]), .B(Key[12]), .Z(n2223) );
  AND2 U2415 ( .A(Key[12]), .B(n2224), .Z(n2219) );
  OR2 U2416 ( .A(n2225), .B(n1974), .Z(n2224) );
  BIC2 U2417 ( .A(n2221), .B(n1975), .Z(n2225) );
  NOT1 U2418 ( .A(Key[76]), .Z(n2221) );
  XOR2 U2419 ( .A(n2226), .B(StateRegOutput[11]), .Z(
        AddKeyConstXOR_XORInst_2_3_N0 ) );
  ORN2 U2420 ( .A(n2227), .B(n2228), .Z(n2226) );
  ORN2 U2421 ( .A(n2229), .B(Key[75]), .Z(n2228) );
  AND2 U2422 ( .A(n2230), .B(n1978), .Z(n2229) );
  OR2 U2423 ( .A(Key[11]), .B(n1975), .Z(n2230) );
  AND2 U2424 ( .A(n2231), .B(Key[11]), .Z(n2227) );
  OR2 U2425 ( .A(n2232), .B(n1974), .Z(n2231) );
  BIC2 U2426 ( .A(n1979), .B(Key[75]), .Z(n2232) );
  XOR2 U2427 ( .A(n2233), .B(StateRegOutput[10]), .Z(
        AddKeyConstXOR_XORInst_2_2_N0 ) );
  ORN2 U2428 ( .A(n2234), .B(n2235), .Z(n2233) );
  ORN2 U2429 ( .A(n2236), .B(Key[74]), .Z(n2235) );
  AND2 U2430 ( .A(n2237), .B(n1978), .Z(n2236) );
  OR2 U2431 ( .A(Key[10]), .B(n1975), .Z(n2237) );
  AND2 U2432 ( .A(n2238), .B(Key[10]), .Z(n2234) );
  OR2 U2433 ( .A(n2239), .B(n1974), .Z(n2238) );
  BIC2 U2434 ( .A(n1979), .B(Key[74]), .Z(n2239) );
  XOR2 U2435 ( .A(n2240), .B(StateRegOutput[9]), .Z(
        AddKeyConstXOR_XORInst_2_1_N0 ) );
  ORN2 U2436 ( .A(n2241), .B(n2242), .Z(n2240) );
  ORN2 U2437 ( .A(n2243), .B(Key[9]), .Z(n2242) );
  BIC2 U2438 ( .A(n2244), .B(n1974), .Z(n2243) );
  OR2 U2439 ( .A(Key[73]), .B(n1975), .Z(n2244) );
  AND2 U2440 ( .A(n2245), .B(Key[73]), .Z(n2241) );
  ORN2 U2441 ( .A(n2246), .B(n1978), .Z(n2245) );
  BIC2 U2442 ( .A(n1979), .B(Key[9]), .Z(n2246) );
  NOT1 U2443 ( .A(n1850), .Z(AddKeyConstXOR_XORInst_2_0_N1 ) );
  XOR2 U2444 ( .A(n2247), .B(n2248), .Z(n1850) );
  AND2 U2445 ( .A(n2249), .B(n1998), .Z(n2248) );
  NOT1 U2446 ( .A(n2250), .Z(n1998) );
  BIC2 U2447 ( .A(n1943), .B(n1953), .Z(n2249) );
  XOR2 U2448 ( .A(n2251), .B(StateRegOutput[8]), .Z(n2247) );
  ORN2 U2449 ( .A(n2252), .B(n2253), .Z(n2251) );
  ORN2 U2450 ( .A(n2254), .B(n2255), .Z(n2253) );
  AND2 U2451 ( .A(n2256), .B(n2005), .Z(n2255) );
  ORN2 U2452 ( .A(n1974), .B(Key[72]), .Z(n2256) );
  AND2 U2453 ( .A(Key[72]), .B(n2257), .Z(n2252) );
  ORN2 U2454 ( .A(n2258), .B(n1978), .Z(n2257) );
  BIC2 U2455 ( .A(n2254), .B(n1975), .Z(n2258) );
  NOT1 U2456 ( .A(Key[8]), .Z(n2254) );
  XOR2 U2457 ( .A(n2259), .B(StateRegOutput[7]), .Z(
        AddKeyConstXOR_XORInst_1_3_N0 ) );
  ORN2 U2458 ( .A(n2260), .B(n2261), .Z(n2259) );
  ORN2 U2459 ( .A(n2262), .B(Key[7]), .Z(n2261) );
  BIC2 U2460 ( .A(n2263), .B(n1974), .Z(n2262) );
  OR2 U2461 ( .A(Key[71]), .B(n1975), .Z(n2263) );
  AND2 U2462 ( .A(n2264), .B(Key[71]), .Z(n2260) );
  ORN2 U2463 ( .A(n2265), .B(n1978), .Z(n2264) );
  BIC2 U2464 ( .A(n1979), .B(Key[7]), .Z(n2265) );
  XOR2 U2465 ( .A(n2266), .B(StateRegOutput[6]), .Z(
        AddKeyConstXOR_XORInst_1_2_N0 ) );
  ORN2 U2466 ( .A(n2267), .B(n2268), .Z(n2266) );
  ORN2 U2467 ( .A(n2269), .B(Key[70]), .Z(n2268) );
  AND2 U2468 ( .A(n2270), .B(n1978), .Z(n2269) );
  OR2 U2469 ( .A(Key[6]), .B(n1975), .Z(n2270) );
  AND2 U2470 ( .A(n2271), .B(Key[6]), .Z(n2267) );
  OR2 U2471 ( .A(n2272), .B(n1974), .Z(n2271) );
  BIC2 U2472 ( .A(n1979), .B(Key[70]), .Z(n2272) );
  XOR2 U2473 ( .A(n2273), .B(StateRegOutput[5]), .Z(
        AddKeyConstXOR_XORInst_1_1_N0 ) );
  ORN2 U2474 ( .A(n2274), .B(n2275), .Z(n2273) );
  ORN2 U2475 ( .A(n2276), .B(Key[69]), .Z(n2275) );
  AND2 U2476 ( .A(n2277), .B(n1978), .Z(n2276) );
  OR2 U2477 ( .A(Key[5]), .B(n1975), .Z(n2277) );
  AND2 U2478 ( .A(n2278), .B(Key[5]), .Z(n2274) );
  OR2 U2479 ( .A(n2279), .B(n1974), .Z(n2278) );
  BIC2 U2480 ( .A(n1979), .B(Key[69]), .Z(n2279) );
  NOT1 U2481 ( .A(n1589), .Z(AddKeyConstXOR_XORInst_1_0_N1 ) );
  XOR2 U2482 ( .A(n2280), .B(n2281), .Z(n1589) );
  AND2 U2483 ( .A(n2282), .B(n2283), .Z(n2281) );
  AND2 U2484 ( .A(n2284), .B(n1943), .Z(n2283) );
  NOT1 U2485 ( .A(n2217), .Z(n1943) );
  AND2 U2486 ( .A(n1946), .B(n2036), .Z(n2217) );
  ORN2 U2487 ( .A(n2036), .B(n1953), .Z(n2284) );
  AND2 U2488 ( .A(n2285), .B(n2286), .Z(n2282) );
  ORN2 U2489 ( .A(n2287), .B(Round[0]), .Z(n2286) );
  XOR2 U2490 ( .A(n2288), .B(StateRegOutput[4]), .Z(n2280) );
  ORN2 U2491 ( .A(n2289), .B(n2290), .Z(n2288) );
  ORN2 U2492 ( .A(n2291), .B(n2292), .Z(n2290) );
  BIC2 U2493 ( .A(n2293), .B(n1974), .Z(n2292) );
  ORN2 U2494 ( .A(Round[0]), .B(Key[4]), .Z(n2293) );
  AND2 U2495 ( .A(Key[4]), .B(n2294), .Z(n2289) );
  OR2 U2496 ( .A(n2295), .B(n1974), .Z(n2294) );
  BIC2 U2497 ( .A(n2291), .B(n1975), .Z(n2295) );
  NOT1 U2498 ( .A(Key[68]), .Z(n2291) );
  XOR2 U2499 ( .A(n2296), .B(StateRegOutput[63]), .Z(
        AddKeyConstXOR_XORInst_15_3_N0 ) );
  ORN2 U2500 ( .A(n2297), .B(n2298), .Z(n2296) );
  ORN2 U2501 ( .A(n2299), .B(Key[63]), .Z(n2298) );
  BIC2 U2502 ( .A(n2300), .B(n1974), .Z(n2299) );
  OR2 U2503 ( .A(Key[127]), .B(n1975), .Z(n2300) );
  AND2 U2504 ( .A(n2301), .B(Key[127]), .Z(n2297) );
  ORN2 U2505 ( .A(n2302), .B(n1978), .Z(n2301) );
  BIC2 U2506 ( .A(n1979), .B(Key[63]), .Z(n2302) );
  XOR2 U2507 ( .A(n2303), .B(StateRegOutput[62]), .Z(
        AddKeyConstXOR_XORInst_15_2_N0 ) );
  ORN2 U2508 ( .A(n2304), .B(n2305), .Z(n2303) );
  ORN2 U2509 ( .A(n2306), .B(Key[62]), .Z(n2305) );
  BIC2 U2510 ( .A(n2307), .B(n1974), .Z(n2306) );
  OR2 U2511 ( .A(Key[126]), .B(n1975), .Z(n2307) );
  AND2 U2512 ( .A(n2308), .B(Key[126]), .Z(n2304) );
  ORN2 U2513 ( .A(n2309), .B(n1978), .Z(n2308) );
  BIC2 U2514 ( .A(n1979), .B(Key[62]), .Z(n2309) );
  XOR2 U2515 ( .A(n2310), .B(StateRegOutput[61]), .Z(
        AddKeyConstXOR_XORInst_15_1_N0 ) );
  ORN2 U2516 ( .A(n2311), .B(n2312), .Z(n2310) );
  ORN2 U2517 ( .A(n2313), .B(Key[61]), .Z(n2312) );
  BIC2 U2518 ( .A(n2314), .B(n1974), .Z(n2313) );
  OR2 U2519 ( .A(Key[125]), .B(n1975), .Z(n2314) );
  AND2 U2520 ( .A(n2315), .B(Key[125]), .Z(n2311) );
  ORN2 U2521 ( .A(n2316), .B(n1978), .Z(n2315) );
  BIC2 U2522 ( .A(n1979), .B(Key[61]), .Z(n2316) );
  NOT1 U2523 ( .A(n1400), .Z(AddKeyConstXOR_XORInst_15_0_N1 ) );
  XOR2 U2524 ( .A(n2317), .B(n2318), .Z(n1400) );
  AND2 U2525 ( .A(n2319), .B(n2320), .Z(n2318) );
  ORN2 U2526 ( .A(n2321), .B(Round[3]), .Z(n2320) );
  AND2 U2527 ( .A(n2322), .B(n2037), .Z(n2321) );
  ORN2 U2528 ( .A(n1964), .B(Round[2]), .Z(n2322) );
  AND2 U2529 ( .A(n2323), .B(n1959), .Z(n2319) );
  NOT1 U2530 ( .A(n1954), .Z(n1959) );
  ORN2 U2531 ( .A(n1964), .B(n2143), .Z(n2323) );
  XOR2 U2532 ( .A(n2324), .B(StateRegOutput[60]), .Z(n2317) );
  ORN2 U2533 ( .A(n2325), .B(n2326), .Z(n2324) );
  ORN2 U2534 ( .A(n2327), .B(n2328), .Z(n2326) );
  AND2 U2535 ( .A(n2329), .B(n2005), .Z(n2328) );
  ORN2 U2536 ( .A(n1974), .B(Key[124]), .Z(n2329) );
  AND2 U2537 ( .A(Key[124]), .B(n2330), .Z(n2325) );
  ORN2 U2538 ( .A(n2331), .B(n1978), .Z(n2330) );
  BIC2 U2539 ( .A(n2327), .B(n1975), .Z(n2331) );
  NOT1 U2540 ( .A(Key[60]), .Z(n2327) );
  XOR2 U2541 ( .A(n2332), .B(StateRegOutput[59]), .Z(
        AddKeyConstXOR_XORInst_14_3_N0 ) );
  ORN2 U2542 ( .A(n2333), .B(n2334), .Z(n2332) );
  ORN2 U2543 ( .A(n2335), .B(Key[59]), .Z(n2334) );
  BIC2 U2544 ( .A(n2336), .B(n1974), .Z(n2335) );
  OR2 U2545 ( .A(Key[123]), .B(n1975), .Z(n2336) );
  AND2 U2546 ( .A(n2337), .B(Key[123]), .Z(n2333) );
  ORN2 U2547 ( .A(n2338), .B(n1978), .Z(n2337) );
  BIC2 U2548 ( .A(n1979), .B(Key[59]), .Z(n2338) );
  XOR2 U2549 ( .A(n2339), .B(StateRegOutput[58]), .Z(
        AddKeyConstXOR_XORInst_14_2_N0 ) );
  ORN2 U2550 ( .A(n2340), .B(n2341), .Z(n2339) );
  ORN2 U2551 ( .A(n2342), .B(Key[58]), .Z(n2341) );
  BIC2 U2552 ( .A(n2343), .B(n1974), .Z(n2342) );
  OR2 U2553 ( .A(Key[122]), .B(n1975), .Z(n2343) );
  AND2 U2554 ( .A(n2344), .B(Key[122]), .Z(n2340) );
  ORN2 U2555 ( .A(n2345), .B(n1978), .Z(n2344) );
  BIC2 U2556 ( .A(n1979), .B(Key[58]), .Z(n2345) );
  XOR2 U2557 ( .A(n2346), .B(StateRegOutput[57]), .Z(
        AddKeyConstXOR_XORInst_14_1_N0 ) );
  ORN2 U2558 ( .A(n2347), .B(n2348), .Z(n2346) );
  ORN2 U2559 ( .A(n2349), .B(Key[57]), .Z(n2348) );
  BIC2 U2560 ( .A(n2350), .B(n1974), .Z(n2349) );
  OR2 U2561 ( .A(Key[121]), .B(n1975), .Z(n2350) );
  AND2 U2562 ( .A(n2351), .B(Key[121]), .Z(n2347) );
  ORN2 U2563 ( .A(n2352), .B(n1978), .Z(n2351) );
  BIC2 U2564 ( .A(n1979), .B(Key[57]), .Z(n2352) );
  NOT1 U2565 ( .A(n1526), .Z(AddKeyConstXOR_XORInst_14_0_N1 ) );
  XOR2 U2566 ( .A(n2353), .B(n2354), .Z(n1526) );
  AND2 U2567 ( .A(n2355), .B(n2356), .Z(n2354) );
  AND2 U2568 ( .A(n2183), .B(n2074), .Z(n2356) );
  NOT1 U2569 ( .A(n2040), .Z(n2074) );
  ORN2 U2570 ( .A(n2357), .B(Round[2]), .Z(n2183) );
  ORN2 U2571 ( .A(Round[0]), .B(n2036), .Z(n2357) );
  AND2 U2572 ( .A(n2358), .B(n2039), .Z(n2355) );
  NOT1 U2573 ( .A(n2149), .Z(n2039) );
  AND2 U2574 ( .A(n1946), .B(Round[3]), .Z(n2149) );
  ORN2 U2575 ( .A(Round[0]), .B(Round[1]), .Z(n2358) );
  XOR2 U2576 ( .A(n2359), .B(StateRegOutput[56]), .Z(n2353) );
  ORN2 U2577 ( .A(n2360), .B(n2361), .Z(n2359) );
  ORN2 U2578 ( .A(n2362), .B(n2363), .Z(n2361) );
  AND2 U2579 ( .A(n2364), .B(n2005), .Z(n2363) );
  ORN2 U2580 ( .A(n1974), .B(Key[120]), .Z(n2364) );
  AND2 U2581 ( .A(Key[120]), .B(n2365), .Z(n2360) );
  ORN2 U2582 ( .A(n2366), .B(n1978), .Z(n2365) );
  BIC2 U2583 ( .A(n2362), .B(n1975), .Z(n2366) );
  NOT1 U2584 ( .A(Key[56]), .Z(n2362) );
  XOR2 U2585 ( .A(n2367), .B(StateRegOutput[55]), .Z(
        AddKeyConstXOR_XORInst_13_3_N0 ) );
  ORN2 U2586 ( .A(n2368), .B(n2369), .Z(n2367) );
  ORN2 U2587 ( .A(n2370), .B(Key[55]), .Z(n2369) );
  BIC2 U2588 ( .A(n2371), .B(n1974), .Z(n2370) );
  OR2 U2589 ( .A(Key[119]), .B(n1975), .Z(n2371) );
  AND2 U2590 ( .A(n2372), .B(Key[119]), .Z(n2368) );
  ORN2 U2591 ( .A(n2373), .B(n1978), .Z(n2372) );
  BIC2 U2592 ( .A(n1979), .B(Key[55]), .Z(n2373) );
  XOR2 U2593 ( .A(n2374), .B(StateRegOutput[54]), .Z(
        AddKeyConstXOR_XORInst_13_2_N0 ) );
  ORN2 U2594 ( .A(n2375), .B(n2376), .Z(n2374) );
  ORN2 U2595 ( .A(n2377), .B(Key[54]), .Z(n2376) );
  BIC2 U2596 ( .A(n2378), .B(n1974), .Z(n2377) );
  OR2 U2597 ( .A(Key[118]), .B(n1975), .Z(n2378) );
  AND2 U2598 ( .A(n2379), .B(Key[118]), .Z(n2375) );
  ORN2 U2599 ( .A(n2380), .B(n1978), .Z(n2379) );
  BIC2 U2600 ( .A(n1979), .B(Key[54]), .Z(n2380) );
  XOR2 U2601 ( .A(n2381), .B(StateRegOutput[53]), .Z(
        AddKeyConstXOR_XORInst_13_1_N0 ) );
  ORN2 U2602 ( .A(n2382), .B(n2383), .Z(n2381) );
  ORN2 U2603 ( .A(n2384), .B(Key[53]), .Z(n2383) );
  BIC2 U2604 ( .A(n2385), .B(n1974), .Z(n2384) );
  OR2 U2605 ( .A(Key[117]), .B(n1975), .Z(n2385) );
  AND2 U2606 ( .A(n2386), .B(Key[117]), .Z(n2382) );
  ORN2 U2607 ( .A(n2387), .B(n1978), .Z(n2386) );
  BIC2 U2608 ( .A(n1979), .B(Key[53]), .Z(n2387) );
  NOT1 U2609 ( .A(n1860), .Z(AddKeyConstXOR_XORInst_13_0_N1 ) );
  XOR2 U2610 ( .A(n2388), .B(n2389), .Z(n1860) );
  AND2 U2611 ( .A(n2390), .B(n2285), .Z(n2389) );
  BIC2 U2612 ( .A(n2391), .B(n2392), .Z(n2285) );
  NOT1 U2613 ( .A(n1955), .Z(n2392) );
  OR2 U2614 ( .A(n2144), .B(n2393), .Z(n1955) );
  ORN2 U2615 ( .A(Round[0]), .B(n1964), .Z(n2393) );
  ORN2 U2616 ( .A(n2144), .B(n2394), .Z(n2391) );
  BIC2 U2617 ( .A(n2395), .B(n1953), .Z(n2390) );
  AND2 U2618 ( .A(n2396), .B(Round[1]), .Z(n1953) );
  ORN2 U2619 ( .A(Round[2]), .B(n2145), .Z(n2395) );
  XOR2 U2620 ( .A(n2397), .B(StateRegOutput[52]), .Z(n2388) );
  ORN2 U2621 ( .A(n2398), .B(n2399), .Z(n2397) );
  ORN2 U2622 ( .A(n2400), .B(n2401), .Z(n2399) );
  AND2 U2623 ( .A(n2402), .B(n2005), .Z(n2401) );
  ORN2 U2624 ( .A(n1974), .B(Key[116]), .Z(n2402) );
  AND2 U2625 ( .A(Key[116]), .B(n2403), .Z(n2398) );
  ORN2 U2626 ( .A(n2404), .B(n1978), .Z(n2403) );
  BIC2 U2627 ( .A(n2400), .B(n1975), .Z(n2404) );
  NOT1 U2628 ( .A(Key[52]), .Z(n2400) );
  XOR2 U2629 ( .A(n2405), .B(StateRegOutput[51]), .Z(
        AddKeyConstXOR_XORInst_12_3_N0 ) );
  ORN2 U2630 ( .A(n2406), .B(n2407), .Z(n2405) );
  ORN2 U2631 ( .A(n2408), .B(Key[51]), .Z(n2407) );
  BIC2 U2632 ( .A(n2409), .B(n1974), .Z(n2408) );
  OR2 U2633 ( .A(Key[115]), .B(n1975), .Z(n2409) );
  AND2 U2634 ( .A(n2410), .B(Key[115]), .Z(n2406) );
  ORN2 U2635 ( .A(n2411), .B(n1978), .Z(n2410) );
  BIC2 U2636 ( .A(n1979), .B(Key[51]), .Z(n2411) );
  XOR2 U2637 ( .A(n2412), .B(StateRegOutput[50]), .Z(
        AddKeyConstXOR_XORInst_12_2_N0 ) );
  ORN2 U2638 ( .A(n2413), .B(n2414), .Z(n2412) );
  ORN2 U2639 ( .A(n2415), .B(Key[50]), .Z(n2414) );
  BIC2 U2640 ( .A(n2416), .B(n1974), .Z(n2415) );
  OR2 U2641 ( .A(Key[114]), .B(n1975), .Z(n2416) );
  AND2 U2642 ( .A(n2417), .B(Key[114]), .Z(n2413) );
  ORN2 U2643 ( .A(n2418), .B(n1978), .Z(n2417) );
  BIC2 U2644 ( .A(n1979), .B(Key[50]), .Z(n2418) );
  XOR2 U2645 ( .A(n2419), .B(StateRegOutput[49]), .Z(
        AddKeyConstXOR_XORInst_12_1_N0 ) );
  ORN2 U2646 ( .A(n2420), .B(n2421), .Z(n2419) );
  ORN2 U2647 ( .A(n2422), .B(Key[49]), .Z(n2421) );
  BIC2 U2648 ( .A(n2423), .B(n1974), .Z(n2422) );
  OR2 U2649 ( .A(Key[113]), .B(n1975), .Z(n2423) );
  AND2 U2650 ( .A(n2424), .B(Key[113]), .Z(n2420) );
  ORN2 U2651 ( .A(n2425), .B(n1978), .Z(n2424) );
  BIC2 U2652 ( .A(n1979), .B(Key[49]), .Z(n2425) );
  NOT1 U2653 ( .A(n1778), .Z(AddKeyConstXOR_XORInst_12_0_N1 ) );
  XOR2 U2654 ( .A(n2426), .B(n2427), .Z(n1778) );
  AND2 U2655 ( .A(n2108), .B(n2428), .Z(n2427) );
  ORN2 U2656 ( .A(n2145), .B(Round[0]), .Z(n2428) );
  BIC2 U2657 ( .A(n2429), .B(n1954), .Z(n2108) );
  AND2 U2658 ( .A(n2430), .B(Round[2]), .Z(n1954) );
  BIC2 U2659 ( .A(Round[1]), .B(Round[0]), .Z(n2430) );
  ORN2 U2660 ( .A(Round[0]), .B(n2145), .Z(n2429) );
  BIC2 U2661 ( .A(n2036), .B(n1964), .Z(n2145) );
  XOR2 U2662 ( .A(n2431), .B(StateRegOutput[48]), .Z(n2426) );
  ORN2 U2663 ( .A(n2432), .B(n2433), .Z(n2431) );
  ORN2 U2664 ( .A(n2434), .B(n2435), .Z(n2433) );
  AND2 U2665 ( .A(n2436), .B(n2005), .Z(n2435) );
  ORN2 U2666 ( .A(n1974), .B(Key[112]), .Z(n2436) );
  AND2 U2667 ( .A(Key[112]), .B(n2437), .Z(n2432) );
  ORN2 U2668 ( .A(n2438), .B(n1978), .Z(n2437) );
  BIC2 U2669 ( .A(n2434), .B(n1975), .Z(n2438) );
  NOT1 U2670 ( .A(Key[48]), .Z(n2434) );
  XOR2 U2671 ( .A(n2439), .B(StateRegOutput[47]), .Z(
        AddKeyConstXOR_XORInst_11_3_N0 ) );
  ORN2 U2672 ( .A(n2440), .B(n2441), .Z(n2439) );
  ORN2 U2673 ( .A(n2442), .B(Key[47]), .Z(n2441) );
  BIC2 U2674 ( .A(n2443), .B(n1974), .Z(n2442) );
  OR2 U2675 ( .A(Key[111]), .B(n1975), .Z(n2443) );
  AND2 U2676 ( .A(n2444), .B(Key[111]), .Z(n2440) );
  ORN2 U2677 ( .A(n2445), .B(n1978), .Z(n2444) );
  BIC2 U2678 ( .A(n1979), .B(Key[47]), .Z(n2445) );
  XOR2 U2679 ( .A(n2446), .B(StateRegOutput[46]), .Z(
        AddKeyConstXOR_XORInst_11_2_N0 ) );
  ORN2 U2680 ( .A(n2447), .B(n2448), .Z(n2446) );
  ORN2 U2681 ( .A(n2449), .B(Key[46]), .Z(n2448) );
  BIC2 U2682 ( .A(n2450), .B(n1974), .Z(n2449) );
  OR2 U2683 ( .A(Key[110]), .B(n1975), .Z(n2450) );
  AND2 U2684 ( .A(n2451), .B(Key[110]), .Z(n2447) );
  ORN2 U2685 ( .A(n2452), .B(n1978), .Z(n2451) );
  BIC2 U2686 ( .A(n1979), .B(Key[46]), .Z(n2452) );
  XOR2 U2687 ( .A(n2453), .B(StateRegOutput[45]), .Z(
        AddKeyConstXOR_XORInst_11_1_N0 ) );
  ORN2 U2688 ( .A(n2454), .B(n2455), .Z(n2453) );
  ORN2 U2689 ( .A(n2456), .B(Key[45]), .Z(n2455) );
  BIC2 U2690 ( .A(n2457), .B(n1974), .Z(n2456) );
  OR2 U2691 ( .A(Key[109]), .B(n1975), .Z(n2457) );
  AND2 U2692 ( .A(n2458), .B(Key[109]), .Z(n2454) );
  ORN2 U2693 ( .A(n2459), .B(n1978), .Z(n2458) );
  BIC2 U2694 ( .A(n1979), .B(Key[45]), .Z(n2459) );
  NOT1 U2695 ( .A(n1581), .Z(AddKeyConstXOR_XORInst_11_0_N1 ) );
  XOR2 U2696 ( .A(n2460), .B(n2461), .Z(n1581) );
  AND2 U2697 ( .A(n2462), .B(n2463), .Z(n2461) );
  ORN2 U2698 ( .A(n2144), .B(n2040), .Z(n2463) );
  AND2 U2699 ( .A(n2464), .B(n2034), .Z(n2462) );
  ORN2 U2700 ( .A(Round[2]), .B(n2250), .Z(n2034) );
  BIC2 U2701 ( .A(n1964), .B(n2075), .Z(n2250) );
  NOT1 U2702 ( .A(n2394), .Z(n2075) );
  BIC2 U2703 ( .A(n1978), .B(n2036), .Z(n2394) );
  ORN2 U2704 ( .A(Round[3]), .B(n2148), .Z(n2464) );
  NOT1 U2705 ( .A(n1960), .Z(n2148) );
  OR2 U2706 ( .A(n1964), .B(n1968), .Z(n1960) );
  XOR2 U2707 ( .A(n2465), .B(StateRegOutput[44]), .Z(n2460) );
  ORN2 U2708 ( .A(n2466), .B(n2467), .Z(n2465) );
  ORN2 U2709 ( .A(n2468), .B(n2469), .Z(n2467) );
  AND2 U2710 ( .A(n2470), .B(n2005), .Z(n2469) );
  ORN2 U2711 ( .A(n1974), .B(Key[108]), .Z(n2470) );
  AND2 U2712 ( .A(Key[108]), .B(n2471), .Z(n2466) );
  ORN2 U2713 ( .A(n2472), .B(n1978), .Z(n2471) );
  BIC2 U2714 ( .A(n2468), .B(n1975), .Z(n2472) );
  NOT1 U2715 ( .A(Key[44]), .Z(n2468) );
  XOR2 U2716 ( .A(n2473), .B(StateRegOutput[43]), .Z(
        AddKeyConstXOR_XORInst_10_3_N0 ) );
  ORN2 U2717 ( .A(n2474), .B(n2475), .Z(n2473) );
  ORN2 U2718 ( .A(n2476), .B(Key[43]), .Z(n2475) );
  BIC2 U2719 ( .A(n2477), .B(n1974), .Z(n2476) );
  OR2 U2720 ( .A(Key[107]), .B(n1975), .Z(n2477) );
  AND2 U2721 ( .A(n2478), .B(Key[107]), .Z(n2474) );
  ORN2 U2722 ( .A(n2479), .B(n1978), .Z(n2478) );
  BIC2 U2723 ( .A(n1979), .B(Key[43]), .Z(n2479) );
  XOR2 U2724 ( .A(n2480), .B(StateRegOutput[42]), .Z(
        AddKeyConstXOR_XORInst_10_2_N0 ) );
  ORN2 U2725 ( .A(n2481), .B(n2482), .Z(n2480) );
  ORN2 U2726 ( .A(n2483), .B(Key[42]), .Z(n2482) );
  BIC2 U2727 ( .A(n2484), .B(n1974), .Z(n2483) );
  OR2 U2728 ( .A(Key[106]), .B(n1975), .Z(n2484) );
  AND2 U2729 ( .A(n2485), .B(Key[106]), .Z(n2481) );
  ORN2 U2730 ( .A(n2486), .B(n1978), .Z(n2485) );
  BIC2 U2731 ( .A(n1979), .B(Key[42]), .Z(n2486) );
  XOR2 U2732 ( .A(n2487), .B(StateRegOutput[41]), .Z(
        AddKeyConstXOR_XORInst_10_1_N0 ) );
  ORN2 U2733 ( .A(n2488), .B(n2489), .Z(n2487) );
  ORN2 U2734 ( .A(n2490), .B(Key[41]), .Z(n2489) );
  BIC2 U2735 ( .A(n2491), .B(n1974), .Z(n2490) );
  OR2 U2736 ( .A(Key[105]), .B(n1975), .Z(n2491) );
  AND2 U2737 ( .A(n2492), .B(Key[105]), .Z(n2488) );
  ORN2 U2738 ( .A(n2493), .B(n1978), .Z(n2492) );
  BIC2 U2739 ( .A(n1979), .B(Key[41]), .Z(n2493) );
  NOT1 U2740 ( .A(n1480), .Z(AddKeyConstXOR_XORInst_10_0_N1 ) );
  XOR2 U2741 ( .A(n2494), .B(n2495), .Z(n1480) );
  BIC2 U2742 ( .A(n2496), .B(n1933), .Z(n2495) );
  AND2 U2743 ( .A(n1946), .B(n2040), .Z(n1933) );
  BIC2 U2744 ( .A(Round[1]), .B(n2036), .Z(n2040) );
  AND2 U2745 ( .A(Round[2]), .B(Round[0]), .Z(n1946) );
  BIC2 U2746 ( .A(n2037), .B(n2143), .Z(n2496) );
  AND2 U2747 ( .A(n2396), .B(n2036), .Z(n2143) );
  NOT1 U2748 ( .A(Round[3]), .Z(n2036) );
  ORN2 U2749 ( .A(Round[1]), .B(n2396), .Z(n2037) );
  XOR2 U2750 ( .A(n2497), .B(StateRegOutput[40]), .Z(n2494) );
  ORN2 U2751 ( .A(n2498), .B(n2499), .Z(n2497) );
  ORN2 U2752 ( .A(n2500), .B(n2501), .Z(n2499) );
  AND2 U2753 ( .A(n2502), .B(n2005), .Z(n2501) );
  OR2 U2754 ( .A(n1974), .B(n1979), .Z(n2005) );
  ORN2 U2755 ( .A(n1974), .B(Key[104]), .Z(n2502) );
  AND2 U2756 ( .A(Key[104]), .B(n2503), .Z(n2498) );
  ORN2 U2757 ( .A(n2504), .B(n1978), .Z(n2503) );
  BIC2 U2758 ( .A(n2500), .B(n1975), .Z(n2504) );
  NOT1 U2759 ( .A(Key[40]), .Z(n2500) );
  XOR2 U2760 ( .A(n2505), .B(StateRegOutput[3]), .Z(
        AddKeyConstXOR_XORInst_0_3_N0 ) );
  ORN2 U2761 ( .A(n2506), .B(n2507), .Z(n2505) );
  ORN2 U2762 ( .A(n2508), .B(Key[67]), .Z(n2507) );
  AND2 U2763 ( .A(n2509), .B(n1978), .Z(n2508) );
  OR2 U2764 ( .A(Key[3]), .B(n1975), .Z(n2509) );
  AND2 U2765 ( .A(n2510), .B(Key[3]), .Z(n2506) );
  OR2 U2766 ( .A(n2511), .B(n1974), .Z(n2510) );
  BIC2 U2767 ( .A(n1979), .B(Key[67]), .Z(n2511) );
  XOR2 U2768 ( .A(n2512), .B(StateRegOutput[2]), .Z(
        AddKeyConstXOR_XORInst_0_2_N0 ) );
  ORN2 U2769 ( .A(n2513), .B(n2514), .Z(n2512) );
  ORN2 U2770 ( .A(n2515), .B(Key[66]), .Z(n2514) );
  AND2 U2771 ( .A(n2516), .B(n1978), .Z(n2515) );
  OR2 U2772 ( .A(Key[2]), .B(n1975), .Z(n2516) );
  AND2 U2773 ( .A(n2517), .B(Key[2]), .Z(n2513) );
  OR2 U2774 ( .A(n2518), .B(n1974), .Z(n2517) );
  BIC2 U2775 ( .A(n1979), .B(Key[66]), .Z(n2518) );
  XOR2 U2776 ( .A(n2519), .B(StateRegOutput[1]), .Z(
        AddKeyConstXOR_XORInst_0_1_N0 ) );
  ORN2 U2777 ( .A(n2520), .B(n2521), .Z(n2519) );
  ORN2 U2778 ( .A(n2522), .B(Key[65]), .Z(n2521) );
  AND2 U2779 ( .A(n2523), .B(n1978), .Z(n2522) );
  OR2 U2780 ( .A(Key[1]), .B(n1975), .Z(n2523) );
  AND2 U2781 ( .A(n2524), .B(Key[1]), .Z(n2520) );
  OR2 U2782 ( .A(n2525), .B(n1974), .Z(n2524) );
  BIC2 U2783 ( .A(n1979), .B(Key[65]), .Z(n2525) );
  NOT1 U2784 ( .A(n1975), .Z(n1979) );
  NOT1 U2785 ( .A(n1517), .Z(AddKeyConstXOR_XORInst_0_0_N1 ) );
  XOR2 U2786 ( .A(n2526), .B(n2527), .Z(n1517) );
  BIC2 U2787 ( .A(n2528), .B(n2396), .Z(n2527) );
  BIC2 U2788 ( .A(n2144), .B(n1978), .Z(n2396) );
  ORN2 U2789 ( .A(n2287), .B(Round[2]), .Z(n2528) );
  XOR2 U2790 ( .A(n2529), .B(StateRegOutput[0]), .Z(n2526) );
  ORN2 U2791 ( .A(n2530), .B(n2531), .Z(n2529) );
  ORN2 U2792 ( .A(n2532), .B(n2533), .Z(n2531) );
  BIC2 U2793 ( .A(n2534), .B(n1974), .Z(n2533) );
  ORN2 U2794 ( .A(Round[0]), .B(Key[0]), .Z(n2534) );
  AND2 U2795 ( .A(Key[0]), .B(n2535), .Z(n2530) );
  OR2 U2796 ( .A(n2536), .B(n1974), .Z(n2535) );
  AND2 U2797 ( .A(n1975), .B(n1978), .Z(n1974) );
  NOT1 U2798 ( .A(Round[0]), .Z(n1978) );
  BIC2 U2799 ( .A(n2532), .B(n1975), .Z(n2536) );
  OR2 U2800 ( .A(n2287), .B(n1968), .Z(n1975) );
  ORN2 U2801 ( .A(Round[0]), .B(n2144), .Z(n1968) );
  NOT1 U2802 ( .A(Round[2]), .Z(n2144) );
  ORN2 U2803 ( .A(Round[3]), .B(n1964), .Z(n2287) );
  NOT1 U2804 ( .A(Round[1]), .Z(n1964) );
  NOT1 U2805 ( .A(Key[64]), .Z(n2532) );
endmodule

