
module LED64Enc ( clk, rst, Plaintext, Key, Ciphertext, done );
  input [63:0] Plaintext;
  input [63:0] Key;
  output [63:0] Ciphertext;
  input clk, rst;
  output done;
  wire   AddKey, PlaintextMUX_MUXInst_0_n2 , PlaintextMUX_MUXInst_0_n1 ,
         PlaintextMUX_MUXInst_1_n2 , PlaintextMUX_MUXInst_1_n1 ,
         PlaintextMUX_MUXInst_2_n2 , PlaintextMUX_MUXInst_2_n1 ,
         PlaintextMUX_MUXInst_3_n2 , PlaintextMUX_MUXInst_3_n1 ,
         PlaintextMUX_MUXInst_4_n2 , PlaintextMUX_MUXInst_4_n1 ,
         PlaintextMUX_MUXInst_5_n2 , PlaintextMUX_MUXInst_5_n1 ,
         PlaintextMUX_MUXInst_6_n2 , PlaintextMUX_MUXInst_6_n1 ,
         PlaintextMUX_MUXInst_7_n2 , PlaintextMUX_MUXInst_7_n1 ,
         PlaintextMUX_MUXInst_8_n2 , PlaintextMUX_MUXInst_8_n1 ,
         PlaintextMUX_MUXInst_9_n2 , PlaintextMUX_MUXInst_9_n1 ,
         PlaintextMUX_MUXInst_10_n2 , PlaintextMUX_MUXInst_10_n1 ,
         PlaintextMUX_MUXInst_11_n2 , PlaintextMUX_MUXInst_11_n1 ,
         PlaintextMUX_MUXInst_12_n2 , PlaintextMUX_MUXInst_12_n1 ,
         PlaintextMUX_MUXInst_13_n2 , PlaintextMUX_MUXInst_13_n1 ,
         PlaintextMUX_MUXInst_14_n2 , PlaintextMUX_MUXInst_14_n1 ,
         PlaintextMUX_MUXInst_15_n2 , PlaintextMUX_MUXInst_15_n1 ,
         PlaintextMUX_MUXInst_16_n2 , PlaintextMUX_MUXInst_16_n1 ,
         PlaintextMUX_MUXInst_17_n2 , PlaintextMUX_MUXInst_17_n1 ,
         PlaintextMUX_MUXInst_18_n2 , PlaintextMUX_MUXInst_18_n1 ,
         PlaintextMUX_MUXInst_19_n2 , PlaintextMUX_MUXInst_19_n1 ,
         PlaintextMUX_MUXInst_20_n2 , PlaintextMUX_MUXInst_20_n1 ,
         PlaintextMUX_MUXInst_21_n2 , PlaintextMUX_MUXInst_21_n1 ,
         PlaintextMUX_MUXInst_22_n2 , PlaintextMUX_MUXInst_22_n1 ,
         PlaintextMUX_MUXInst_23_n2 , PlaintextMUX_MUXInst_23_n1 ,
         PlaintextMUX_MUXInst_24_n2 , PlaintextMUX_MUXInst_24_n1 ,
         PlaintextMUX_MUXInst_25_n2 , PlaintextMUX_MUXInst_25_n1 ,
         PlaintextMUX_MUXInst_26_n2 , PlaintextMUX_MUXInst_26_n1 ,
         PlaintextMUX_MUXInst_27_n2 , PlaintextMUX_MUXInst_27_n1 ,
         PlaintextMUX_MUXInst_28_n2 , PlaintextMUX_MUXInst_28_n1 ,
         PlaintextMUX_MUXInst_29_n2 , PlaintextMUX_MUXInst_29_n1 ,
         PlaintextMUX_MUXInst_30_n2 , PlaintextMUX_MUXInst_30_n1 ,
         PlaintextMUX_MUXInst_31_n2 , PlaintextMUX_MUXInst_31_n1 ,
         PlaintextMUX_MUXInst_32_n2 , PlaintextMUX_MUXInst_32_n1 ,
         PlaintextMUX_MUXInst_33_n2 , PlaintextMUX_MUXInst_33_n1 ,
         PlaintextMUX_MUXInst_34_n2 , PlaintextMUX_MUXInst_34_n1 ,
         PlaintextMUX_MUXInst_35_n2 , PlaintextMUX_MUXInst_35_n1 ,
         PlaintextMUX_MUXInst_36_n2 , PlaintextMUX_MUXInst_36_n1 ,
         PlaintextMUX_MUXInst_37_n2 , PlaintextMUX_MUXInst_37_n1 ,
         PlaintextMUX_MUXInst_38_n2 , PlaintextMUX_MUXInst_38_n1 ,
         PlaintextMUX_MUXInst_39_n2 , PlaintextMUX_MUXInst_39_n1 ,
         PlaintextMUX_MUXInst_40_n2 , PlaintextMUX_MUXInst_40_n1 ,
         PlaintextMUX_MUXInst_41_n2 , PlaintextMUX_MUXInst_41_n1 ,
         PlaintextMUX_MUXInst_42_n2 , PlaintextMUX_MUXInst_42_n1 ,
         PlaintextMUX_MUXInst_43_n2 , PlaintextMUX_MUXInst_43_n1 ,
         PlaintextMUX_MUXInst_44_n2 , PlaintextMUX_MUXInst_44_n1 ,
         PlaintextMUX_MUXInst_45_n2 , PlaintextMUX_MUXInst_45_n1 ,
         PlaintextMUX_MUXInst_46_n2 , PlaintextMUX_MUXInst_46_n1 ,
         PlaintextMUX_MUXInst_47_n2 , PlaintextMUX_MUXInst_47_n1 ,
         PlaintextMUX_MUXInst_48_n2 , PlaintextMUX_MUXInst_48_n1 ,
         PlaintextMUX_MUXInst_49_n2 , PlaintextMUX_MUXInst_49_n1 ,
         PlaintextMUX_MUXInst_50_n2 , PlaintextMUX_MUXInst_50_n1 ,
         PlaintextMUX_MUXInst_51_n2 , PlaintextMUX_MUXInst_51_n1 ,
         PlaintextMUX_MUXInst_52_n2 , PlaintextMUX_MUXInst_52_n1 ,
         PlaintextMUX_MUXInst_53_n2 , PlaintextMUX_MUXInst_53_n1 ,
         PlaintextMUX_MUXInst_54_n2 , PlaintextMUX_MUXInst_54_n1 ,
         PlaintextMUX_MUXInst_55_n2 , PlaintextMUX_MUXInst_55_n1 ,
         PlaintextMUX_MUXInst_56_n2 , PlaintextMUX_MUXInst_56_n1 ,
         PlaintextMUX_MUXInst_57_n2 , PlaintextMUX_MUXInst_57_n1 ,
         PlaintextMUX_MUXInst_58_n2 , PlaintextMUX_MUXInst_58_n1 ,
         PlaintextMUX_MUXInst_59_n2 , PlaintextMUX_MUXInst_59_n1 ,
         PlaintextMUX_MUXInst_60_n2 , PlaintextMUX_MUXInst_60_n1 ,
         PlaintextMUX_MUXInst_61_n2 , PlaintextMUX_MUXInst_61_n1 ,
         PlaintextMUX_MUXInst_62_n2 , PlaintextMUX_MUXInst_62_n1 ,
         PlaintextMUX_MUXInst_63_n2 , PlaintextMUX_MUXInst_63_n1 ,
         AddKeyXOR_XORInst_0_0_n1 , AddKeyXOR_XORInst_0_1_n1 ,
         AddKeyXOR_XORInst_0_2_n1 , AddKeyXOR_XORInst_0_3_n1 ,
         AddKeyXOR_XORInst_1_0_n1 , AddKeyXOR_XORInst_1_1_n1 ,
         AddKeyXOR_XORInst_1_2_n1 , AddKeyXOR_XORInst_1_3_n1 ,
         AddKeyXOR_XORInst_2_0_n1 , AddKeyXOR_XORInst_2_1_n1 ,
         AddKeyXOR_XORInst_2_2_n1 , AddKeyXOR_XORInst_2_3_n1 ,
         AddKeyXOR_XORInst_3_0_n1 , AddKeyXOR_XORInst_3_1_n1 ,
         AddKeyXOR_XORInst_3_2_n1 , AddKeyXOR_XORInst_3_3_n1 ,
         AddKeyXOR_XORInst_4_0_n1 , AddKeyXOR_XORInst_4_1_n1 ,
         AddKeyXOR_XORInst_4_2_n1 , AddKeyXOR_XORInst_4_3_n1 ,
         AddKeyXOR_XORInst_5_0_n1 , AddKeyXOR_XORInst_5_1_n1 ,
         AddKeyXOR_XORInst_5_2_n1 , AddKeyXOR_XORInst_5_3_n1 ,
         AddKeyXOR_XORInst_6_0_n1 , AddKeyXOR_XORInst_6_1_n1 ,
         AddKeyXOR_XORInst_6_2_n1 , AddKeyXOR_XORInst_6_3_n1 ,
         AddKeyXOR_XORInst_7_0_n1 , AddKeyXOR_XORInst_7_1_n1 ,
         AddKeyXOR_XORInst_7_2_n1 , AddKeyXOR_XORInst_7_3_n1 ,
         AddKeyXOR_XORInst_8_0_n1 , AddKeyXOR_XORInst_8_1_n1 ,
         AddKeyXOR_XORInst_8_2_n1 , AddKeyXOR_XORInst_8_3_n1 ,
         AddKeyXOR_XORInst_9_0_n1 , AddKeyXOR_XORInst_9_1_n1 ,
         AddKeyXOR_XORInst_9_2_n1 , AddKeyXOR_XORInst_9_3_n1 ,
         AddKeyXOR_XORInst_10_0_n1 , AddKeyXOR_XORInst_10_1_n1 ,
         AddKeyXOR_XORInst_10_2_n1 , AddKeyXOR_XORInst_10_3_n1 ,
         AddKeyXOR_XORInst_11_0_n1 , AddKeyXOR_XORInst_11_1_n1 ,
         AddKeyXOR_XORInst_11_2_n1 , AddKeyXOR_XORInst_11_3_n1 ,
         AddKeyXOR_XORInst_12_0_n1 , AddKeyXOR_XORInst_12_1_n1 ,
         AddKeyXOR_XORInst_12_2_n1 , AddKeyXOR_XORInst_12_3_n1 ,
         AddKeyXOR_XORInst_13_0_n1 , AddKeyXOR_XORInst_13_1_n1 ,
         AddKeyXOR_XORInst_13_2_n1 , AddKeyXOR_XORInst_13_3_n1 ,
         AddKeyXOR_XORInst_14_0_n1 , AddKeyXOR_XORInst_14_1_n1 ,
         AddKeyXOR_XORInst_14_2_n1 , AddKeyXOR_XORInst_14_3_n1 ,
         AddKeyXOR_XORInst_15_0_n1 , AddKeyXOR_XORInst_15_1_n1 ,
         AddKeyXOR_XORInst_15_2_n1 , AddKeyXOR_XORInst_15_3_n1 ,
         AddKeyMUX_MUXInst_0_n2 , AddKeyMUX_MUXInst_0_n1 ,
         AddKeyMUX_MUXInst_1_n2 , AddKeyMUX_MUXInst_1_n1 ,
         AddKeyMUX_MUXInst_2_n2 , AddKeyMUX_MUXInst_2_n1 ,
         AddKeyMUX_MUXInst_3_n2 , AddKeyMUX_MUXInst_3_n1 ,
         AddKeyMUX_MUXInst_4_n2 , AddKeyMUX_MUXInst_4_n1 ,
         AddKeyMUX_MUXInst_5_n2 , AddKeyMUX_MUXInst_5_n1 ,
         AddKeyMUX_MUXInst_6_n2 , AddKeyMUX_MUXInst_6_n1 ,
         AddKeyMUX_MUXInst_7_n2 , AddKeyMUX_MUXInst_7_n1 ,
         AddKeyMUX_MUXInst_8_n2 , AddKeyMUX_MUXInst_8_n1 ,
         AddKeyMUX_MUXInst_9_n2 , AddKeyMUX_MUXInst_9_n1 ,
         AddKeyMUX_MUXInst_10_n2 , AddKeyMUX_MUXInst_10_n1 ,
         AddKeyMUX_MUXInst_11_n2 , AddKeyMUX_MUXInst_11_n1 ,
         AddKeyMUX_MUXInst_12_n2 , AddKeyMUX_MUXInst_12_n1 ,
         AddKeyMUX_MUXInst_13_n2 , AddKeyMUX_MUXInst_13_n1 ,
         AddKeyMUX_MUXInst_14_n2 , AddKeyMUX_MUXInst_14_n1 ,
         AddKeyMUX_MUXInst_15_n2 , AddKeyMUX_MUXInst_15_n1 ,
         AddKeyMUX_MUXInst_16_n2 , AddKeyMUX_MUXInst_16_n1 ,
         AddKeyMUX_MUXInst_17_n2 , AddKeyMUX_MUXInst_17_n1 ,
         AddKeyMUX_MUXInst_18_n2 , AddKeyMUX_MUXInst_18_n1 ,
         AddKeyMUX_MUXInst_19_n2 , AddKeyMUX_MUXInst_19_n1 ,
         AddKeyMUX_MUXInst_20_n2 , AddKeyMUX_MUXInst_20_n1 ,
         AddKeyMUX_MUXInst_21_n2 , AddKeyMUX_MUXInst_21_n1 ,
         AddKeyMUX_MUXInst_22_n2 , AddKeyMUX_MUXInst_22_n1 ,
         AddKeyMUX_MUXInst_23_n2 , AddKeyMUX_MUXInst_23_n1 ,
         AddKeyMUX_MUXInst_24_n2 , AddKeyMUX_MUXInst_24_n1 ,
         AddKeyMUX_MUXInst_25_n2 , AddKeyMUX_MUXInst_25_n1 ,
         AddKeyMUX_MUXInst_26_n2 , AddKeyMUX_MUXInst_26_n1 ,
         AddKeyMUX_MUXInst_27_n2 , AddKeyMUX_MUXInst_27_n1 ,
         AddKeyMUX_MUXInst_28_n2 , AddKeyMUX_MUXInst_28_n1 ,
         AddKeyMUX_MUXInst_29_n2 , AddKeyMUX_MUXInst_29_n1 ,
         AddKeyMUX_MUXInst_30_n2 , AddKeyMUX_MUXInst_30_n1 ,
         AddKeyMUX_MUXInst_31_n2 , AddKeyMUX_MUXInst_31_n1 ,
         AddKeyMUX_MUXInst_32_n2 , AddKeyMUX_MUXInst_32_n1 ,
         AddKeyMUX_MUXInst_33_n2 , AddKeyMUX_MUXInst_33_n1 ,
         AddKeyMUX_MUXInst_34_n2 , AddKeyMUX_MUXInst_34_n1 ,
         AddKeyMUX_MUXInst_35_n2 , AddKeyMUX_MUXInst_35_n1 ,
         AddKeyMUX_MUXInst_36_n2 , AddKeyMUX_MUXInst_36_n1 ,
         AddKeyMUX_MUXInst_37_n2 , AddKeyMUX_MUXInst_37_n1 ,
         AddKeyMUX_MUXInst_38_n2 , AddKeyMUX_MUXInst_38_n1 ,
         AddKeyMUX_MUXInst_39_n2 , AddKeyMUX_MUXInst_39_n1 ,
         AddKeyMUX_MUXInst_40_n2 , AddKeyMUX_MUXInst_40_n1 ,
         AddKeyMUX_MUXInst_41_n2 , AddKeyMUX_MUXInst_41_n1 ,
         AddKeyMUX_MUXInst_42_n2 , AddKeyMUX_MUXInst_42_n1 ,
         AddKeyMUX_MUXInst_43_n2 , AddKeyMUX_MUXInst_43_n1 ,
         AddKeyMUX_MUXInst_44_n2 , AddKeyMUX_MUXInst_44_n1 ,
         AddKeyMUX_MUXInst_45_n2 , AddKeyMUX_MUXInst_45_n1 ,
         AddKeyMUX_MUXInst_46_n2 , AddKeyMUX_MUXInst_46_n1 ,
         AddKeyMUX_MUXInst_47_n2 , AddKeyMUX_MUXInst_47_n1 ,
         AddKeyMUX_MUXInst_48_n2 , AddKeyMUX_MUXInst_48_n1 ,
         AddKeyMUX_MUXInst_49_n2 , AddKeyMUX_MUXInst_49_n1 ,
         AddKeyMUX_MUXInst_50_n2 , AddKeyMUX_MUXInst_50_n1 ,
         AddKeyMUX_MUXInst_51_n2 , AddKeyMUX_MUXInst_51_n1 ,
         AddKeyMUX_MUXInst_52_n2 , AddKeyMUX_MUXInst_52_n1 ,
         AddKeyMUX_MUXInst_53_n2 , AddKeyMUX_MUXInst_53_n1 ,
         AddKeyMUX_MUXInst_54_n2 , AddKeyMUX_MUXInst_54_n1 ,
         AddKeyMUX_MUXInst_55_n2 , AddKeyMUX_MUXInst_55_n1 ,
         AddKeyMUX_MUXInst_56_n2 , AddKeyMUX_MUXInst_56_n1 ,
         AddKeyMUX_MUXInst_57_n2 , AddKeyMUX_MUXInst_57_n1 ,
         AddKeyMUX_MUXInst_58_n2 , AddKeyMUX_MUXInst_58_n1 ,
         AddKeyMUX_MUXInst_59_n2 , AddKeyMUX_MUXInst_59_n1 ,
         AddKeyMUX_MUXInst_60_n2 , AddKeyMUX_MUXInst_60_n1 ,
         AddKeyMUX_MUXInst_61_n2 , AddKeyMUX_MUXInst_61_n1 ,
         AddKeyMUX_MUXInst_62_n2 , AddKeyMUX_MUXInst_62_n1 ,
         AddKeyMUX_MUXInst_63_n2 , AddKeyMUX_MUXInst_63_n1 ,
         AddConstXOR_XORInst_XORInst_0_0_n1 ,
         AddConstXOR_XORInst_XORInst_0_1_n1 ,
         AddConstXOR_XORInst_XORInst_0_2_n1 ,
         AddConstXOR_XORInst_XORInst_0_3_n1 ,
         AddConstXOR_XORInst_XORInst_1_0_n1 ,
         AddConstXOR_XORInst_XORInst_1_1_n1 ,
         AddConstXOR_XORInst_XORInst_1_2_n1 ,
         AddConstXOR_XORInst_XORInst_1_3_n1 ,
         AddConstXOR_XORInst_XORInst_2_0_n1 ,
         AddConstXOR_XORInst_XORInst_2_1_n1 ,
         AddConstXOR_XORInst_XORInst_2_2_n1 ,
         AddConstXOR_XORInst_XORInst_2_3_n1 ,
         AddConstXOR_XORInst_XORInst_3_0_n1 ,
         AddConstXOR_XORInst_XORInst_3_1_n1 ,
         AddConstXOR_XORInst_XORInst_3_2_n1 ,
         AddConstXOR_XORInst_XORInst_3_3_n1 ,
         AddConstXOR_XORInst_XORInst_4_0_n1 ,
         AddConstXOR_XORInst_XORInst_4_1_n1 ,
         AddConstXOR_XORInst_XORInst_4_2_n1 ,
         AddConstXOR_XORInst_XORInst_4_3_n1 ,
         AddConstXOR_XORInst_XORInst_5_0_n1 ,
         AddConstXOR_XORInst_XORInst_5_1_n1 ,
         AddConstXOR_XORInst_XORInst_5_2_n1 ,
         AddConstXOR_XORInst_XORInst_5_3_n1 ,
         AddConstXOR_XORInst_XORInst_6_0_n1 ,
         AddConstXOR_XORInst_XORInst_6_1_n1 ,
         AddConstXOR_XORInst_XORInst_6_2_n1 ,
         AddConstXOR_XORInst_XORInst_6_3_n1 ,
         AddConstXOR_XORInst_XORInst_7_0_n1 ,
         AddConstXOR_XORInst_XORInst_7_1_n1 ,
         AddConstXOR_XORInst_XORInst_7_2_n1 ,
         AddConstXOR_XORInst_XORInst_7_3_n1 ,
         SubCellInst_LFInst_0_LFInst_3_n8 ,
         SubCellInst_LFInst_0_LFInst_3_n7 ,
         SubCellInst_LFInst_0_LFInst_3_n6 ,
         SubCellInst_LFInst_0_LFInst_3_n5 ,
         SubCellInst_LFInst_0_LFInst_3_n4 ,
         SubCellInst_LFInst_0_LFInst_3_n3 ,
         SubCellInst_LFInst_0_LFInst_3_n2 ,
         SubCellInst_LFInst_0_LFInst_3_n1 ,
         SubCellInst_LFInst_0_LFInst_2_n10 ,
         SubCellInst_LFInst_0_LFInst_2_n9 ,
         SubCellInst_LFInst_0_LFInst_2_n8 ,
         SubCellInst_LFInst_0_LFInst_2_n7 ,
         SubCellInst_LFInst_0_LFInst_2_n6 ,
         SubCellInst_LFInst_0_LFInst_2_n5 ,
         SubCellInst_LFInst_0_LFInst_2_n4 ,
         SubCellInst_LFInst_0_LFInst_2_n3 ,
         SubCellInst_LFInst_0_LFInst_2_n2 ,
         SubCellInst_LFInst_0_LFInst_2_n1 ,
         SubCellInst_LFInst_0_LFInst_1_n7 ,
         SubCellInst_LFInst_0_LFInst_1_n6 ,
         SubCellInst_LFInst_0_LFInst_1_n5 ,
         SubCellInst_LFInst_0_LFInst_1_n4 ,
         SubCellInst_LFInst_0_LFInst_1_n3 ,
         SubCellInst_LFInst_0_LFInst_1_n2 ,
         SubCellInst_LFInst_0_LFInst_1_n1 ,
         SubCellInst_LFInst_0_LFInst_0_n2 ,
         SubCellInst_LFInst_0_LFInst_0_n1 ,
         SubCellInst_LFInst_1_LFInst_3_n8 ,
         SubCellInst_LFInst_1_LFInst_3_n7 ,
         SubCellInst_LFInst_1_LFInst_3_n6 ,
         SubCellInst_LFInst_1_LFInst_3_n5 ,
         SubCellInst_LFInst_1_LFInst_3_n4 ,
         SubCellInst_LFInst_1_LFInst_3_n3 ,
         SubCellInst_LFInst_1_LFInst_3_n2 ,
         SubCellInst_LFInst_1_LFInst_3_n1 ,
         SubCellInst_LFInst_1_LFInst_2_n10 ,
         SubCellInst_LFInst_1_LFInst_2_n9 ,
         SubCellInst_LFInst_1_LFInst_2_n8 ,
         SubCellInst_LFInst_1_LFInst_2_n7 ,
         SubCellInst_LFInst_1_LFInst_2_n6 ,
         SubCellInst_LFInst_1_LFInst_2_n5 ,
         SubCellInst_LFInst_1_LFInst_2_n4 ,
         SubCellInst_LFInst_1_LFInst_2_n3 ,
         SubCellInst_LFInst_1_LFInst_2_n2 ,
         SubCellInst_LFInst_1_LFInst_2_n1 ,
         SubCellInst_LFInst_1_LFInst_1_n7 ,
         SubCellInst_LFInst_1_LFInst_1_n6 ,
         SubCellInst_LFInst_1_LFInst_1_n5 ,
         SubCellInst_LFInst_1_LFInst_1_n4 ,
         SubCellInst_LFInst_1_LFInst_1_n3 ,
         SubCellInst_LFInst_1_LFInst_1_n2 ,
         SubCellInst_LFInst_1_LFInst_1_n1 ,
         SubCellInst_LFInst_1_LFInst_0_n2 ,
         SubCellInst_LFInst_1_LFInst_0_n1 ,
         SubCellInst_LFInst_2_LFInst_3_n8 ,
         SubCellInst_LFInst_2_LFInst_3_n7 ,
         SubCellInst_LFInst_2_LFInst_3_n6 ,
         SubCellInst_LFInst_2_LFInst_3_n5 ,
         SubCellInst_LFInst_2_LFInst_3_n4 ,
         SubCellInst_LFInst_2_LFInst_3_n3 ,
         SubCellInst_LFInst_2_LFInst_3_n2 ,
         SubCellInst_LFInst_2_LFInst_3_n1 ,
         SubCellInst_LFInst_2_LFInst_2_n10 ,
         SubCellInst_LFInst_2_LFInst_2_n9 ,
         SubCellInst_LFInst_2_LFInst_2_n8 ,
         SubCellInst_LFInst_2_LFInst_2_n7 ,
         SubCellInst_LFInst_2_LFInst_2_n6 ,
         SubCellInst_LFInst_2_LFInst_2_n5 ,
         SubCellInst_LFInst_2_LFInst_2_n4 ,
         SubCellInst_LFInst_2_LFInst_2_n3 ,
         SubCellInst_LFInst_2_LFInst_2_n2 ,
         SubCellInst_LFInst_2_LFInst_2_n1 ,
         SubCellInst_LFInst_2_LFInst_1_n7 ,
         SubCellInst_LFInst_2_LFInst_1_n6 ,
         SubCellInst_LFInst_2_LFInst_1_n5 ,
         SubCellInst_LFInst_2_LFInst_1_n4 ,
         SubCellInst_LFInst_2_LFInst_1_n3 ,
         SubCellInst_LFInst_2_LFInst_1_n2 ,
         SubCellInst_LFInst_2_LFInst_1_n1 ,
         SubCellInst_LFInst_2_LFInst_0_n2 ,
         SubCellInst_LFInst_2_LFInst_0_n1 ,
         SubCellInst_LFInst_3_LFInst_3_n8 ,
         SubCellInst_LFInst_3_LFInst_3_n7 ,
         SubCellInst_LFInst_3_LFInst_3_n6 ,
         SubCellInst_LFInst_3_LFInst_3_n5 ,
         SubCellInst_LFInst_3_LFInst_3_n4 ,
         SubCellInst_LFInst_3_LFInst_3_n3 ,
         SubCellInst_LFInst_3_LFInst_3_n2 ,
         SubCellInst_LFInst_3_LFInst_3_n1 ,
         SubCellInst_LFInst_3_LFInst_2_n10 ,
         SubCellInst_LFInst_3_LFInst_2_n9 ,
         SubCellInst_LFInst_3_LFInst_2_n8 ,
         SubCellInst_LFInst_3_LFInst_2_n7 ,
         SubCellInst_LFInst_3_LFInst_2_n6 ,
         SubCellInst_LFInst_3_LFInst_2_n5 ,
         SubCellInst_LFInst_3_LFInst_2_n4 ,
         SubCellInst_LFInst_3_LFInst_2_n3 ,
         SubCellInst_LFInst_3_LFInst_2_n2 ,
         SubCellInst_LFInst_3_LFInst_2_n1 ,
         SubCellInst_LFInst_3_LFInst_1_n7 ,
         SubCellInst_LFInst_3_LFInst_1_n6 ,
         SubCellInst_LFInst_3_LFInst_1_n5 ,
         SubCellInst_LFInst_3_LFInst_1_n4 ,
         SubCellInst_LFInst_3_LFInst_1_n3 ,
         SubCellInst_LFInst_3_LFInst_1_n2 ,
         SubCellInst_LFInst_3_LFInst_1_n1 ,
         SubCellInst_LFInst_3_LFInst_0_n2 ,
         SubCellInst_LFInst_3_LFInst_0_n1 ,
         SubCellInst_LFInst_4_LFInst_3_n8 ,
         SubCellInst_LFInst_4_LFInst_3_n7 ,
         SubCellInst_LFInst_4_LFInst_3_n6 ,
         SubCellInst_LFInst_4_LFInst_3_n5 ,
         SubCellInst_LFInst_4_LFInst_3_n4 ,
         SubCellInst_LFInst_4_LFInst_3_n3 ,
         SubCellInst_LFInst_4_LFInst_3_n2 ,
         SubCellInst_LFInst_4_LFInst_3_n1 ,
         SubCellInst_LFInst_4_LFInst_2_n10 ,
         SubCellInst_LFInst_4_LFInst_2_n9 ,
         SubCellInst_LFInst_4_LFInst_2_n8 ,
         SubCellInst_LFInst_4_LFInst_2_n7 ,
         SubCellInst_LFInst_4_LFInst_2_n6 ,
         SubCellInst_LFInst_4_LFInst_2_n5 ,
         SubCellInst_LFInst_4_LFInst_2_n4 ,
         SubCellInst_LFInst_4_LFInst_2_n3 ,
         SubCellInst_LFInst_4_LFInst_2_n2 ,
         SubCellInst_LFInst_4_LFInst_2_n1 ,
         SubCellInst_LFInst_4_LFInst_1_n7 ,
         SubCellInst_LFInst_4_LFInst_1_n6 ,
         SubCellInst_LFInst_4_LFInst_1_n5 ,
         SubCellInst_LFInst_4_LFInst_1_n4 ,
         SubCellInst_LFInst_4_LFInst_1_n3 ,
         SubCellInst_LFInst_4_LFInst_1_n2 ,
         SubCellInst_LFInst_4_LFInst_1_n1 ,
         SubCellInst_LFInst_4_LFInst_0_n2 ,
         SubCellInst_LFInst_4_LFInst_0_n1 ,
         SubCellInst_LFInst_5_LFInst_3_n8 ,
         SubCellInst_LFInst_5_LFInst_3_n7 ,
         SubCellInst_LFInst_5_LFInst_3_n6 ,
         SubCellInst_LFInst_5_LFInst_3_n5 ,
         SubCellInst_LFInst_5_LFInst_3_n4 ,
         SubCellInst_LFInst_5_LFInst_3_n3 ,
         SubCellInst_LFInst_5_LFInst_3_n2 ,
         SubCellInst_LFInst_5_LFInst_3_n1 ,
         SubCellInst_LFInst_5_LFInst_2_n10 ,
         SubCellInst_LFInst_5_LFInst_2_n9 ,
         SubCellInst_LFInst_5_LFInst_2_n8 ,
         SubCellInst_LFInst_5_LFInst_2_n7 ,
         SubCellInst_LFInst_5_LFInst_2_n6 ,
         SubCellInst_LFInst_5_LFInst_2_n5 ,
         SubCellInst_LFInst_5_LFInst_2_n4 ,
         SubCellInst_LFInst_5_LFInst_2_n3 ,
         SubCellInst_LFInst_5_LFInst_2_n2 ,
         SubCellInst_LFInst_5_LFInst_2_n1 ,
         SubCellInst_LFInst_5_LFInst_1_n7 ,
         SubCellInst_LFInst_5_LFInst_1_n6 ,
         SubCellInst_LFInst_5_LFInst_1_n5 ,
         SubCellInst_LFInst_5_LFInst_1_n4 ,
         SubCellInst_LFInst_5_LFInst_1_n3 ,
         SubCellInst_LFInst_5_LFInst_1_n2 ,
         SubCellInst_LFInst_5_LFInst_1_n1 ,
         SubCellInst_LFInst_5_LFInst_0_n2 ,
         SubCellInst_LFInst_5_LFInst_0_n1 ,
         SubCellInst_LFInst_6_LFInst_3_n8 ,
         SubCellInst_LFInst_6_LFInst_3_n7 ,
         SubCellInst_LFInst_6_LFInst_3_n6 ,
         SubCellInst_LFInst_6_LFInst_3_n5 ,
         SubCellInst_LFInst_6_LFInst_3_n4 ,
         SubCellInst_LFInst_6_LFInst_3_n3 ,
         SubCellInst_LFInst_6_LFInst_3_n2 ,
         SubCellInst_LFInst_6_LFInst_3_n1 ,
         SubCellInst_LFInst_6_LFInst_2_n10 ,
         SubCellInst_LFInst_6_LFInst_2_n9 ,
         SubCellInst_LFInst_6_LFInst_2_n8 ,
         SubCellInst_LFInst_6_LFInst_2_n7 ,
         SubCellInst_LFInst_6_LFInst_2_n6 ,
         SubCellInst_LFInst_6_LFInst_2_n5 ,
         SubCellInst_LFInst_6_LFInst_2_n4 ,
         SubCellInst_LFInst_6_LFInst_2_n3 ,
         SubCellInst_LFInst_6_LFInst_2_n2 ,
         SubCellInst_LFInst_6_LFInst_2_n1 ,
         SubCellInst_LFInst_6_LFInst_1_n7 ,
         SubCellInst_LFInst_6_LFInst_1_n6 ,
         SubCellInst_LFInst_6_LFInst_1_n5 ,
         SubCellInst_LFInst_6_LFInst_1_n4 ,
         SubCellInst_LFInst_6_LFInst_1_n3 ,
         SubCellInst_LFInst_6_LFInst_1_n2 ,
         SubCellInst_LFInst_6_LFInst_1_n1 ,
         SubCellInst_LFInst_6_LFInst_0_n2 ,
         SubCellInst_LFInst_6_LFInst_0_n1 ,
         SubCellInst_LFInst_7_LFInst_3_n8 ,
         SubCellInst_LFInst_7_LFInst_3_n7 ,
         SubCellInst_LFInst_7_LFInst_3_n6 ,
         SubCellInst_LFInst_7_LFInst_3_n5 ,
         SubCellInst_LFInst_7_LFInst_3_n4 ,
         SubCellInst_LFInst_7_LFInst_3_n3 ,
         SubCellInst_LFInst_7_LFInst_3_n2 ,
         SubCellInst_LFInst_7_LFInst_3_n1 ,
         SubCellInst_LFInst_7_LFInst_2_n10 ,
         SubCellInst_LFInst_7_LFInst_2_n9 ,
         SubCellInst_LFInst_7_LFInst_2_n8 ,
         SubCellInst_LFInst_7_LFInst_2_n7 ,
         SubCellInst_LFInst_7_LFInst_2_n6 ,
         SubCellInst_LFInst_7_LFInst_2_n5 ,
         SubCellInst_LFInst_7_LFInst_2_n4 ,
         SubCellInst_LFInst_7_LFInst_2_n3 ,
         SubCellInst_LFInst_7_LFInst_2_n2 ,
         SubCellInst_LFInst_7_LFInst_2_n1 ,
         SubCellInst_LFInst_7_LFInst_1_n7 ,
         SubCellInst_LFInst_7_LFInst_1_n6 ,
         SubCellInst_LFInst_7_LFInst_1_n5 ,
         SubCellInst_LFInst_7_LFInst_1_n4 ,
         SubCellInst_LFInst_7_LFInst_1_n3 ,
         SubCellInst_LFInst_7_LFInst_1_n2 ,
         SubCellInst_LFInst_7_LFInst_1_n1 ,
         SubCellInst_LFInst_7_LFInst_0_n2 ,
         SubCellInst_LFInst_7_LFInst_0_n1 ,
         SubCellInst_LFInst_8_LFInst_3_n8 ,
         SubCellInst_LFInst_8_LFInst_3_n7 ,
         SubCellInst_LFInst_8_LFInst_3_n6 ,
         SubCellInst_LFInst_8_LFInst_3_n5 ,
         SubCellInst_LFInst_8_LFInst_3_n4 ,
         SubCellInst_LFInst_8_LFInst_3_n3 ,
         SubCellInst_LFInst_8_LFInst_3_n2 ,
         SubCellInst_LFInst_8_LFInst_3_n1 ,
         SubCellInst_LFInst_8_LFInst_2_n10 ,
         SubCellInst_LFInst_8_LFInst_2_n9 ,
         SubCellInst_LFInst_8_LFInst_2_n8 ,
         SubCellInst_LFInst_8_LFInst_2_n7 ,
         SubCellInst_LFInst_8_LFInst_2_n6 ,
         SubCellInst_LFInst_8_LFInst_2_n5 ,
         SubCellInst_LFInst_8_LFInst_2_n4 ,
         SubCellInst_LFInst_8_LFInst_2_n3 ,
         SubCellInst_LFInst_8_LFInst_2_n2 ,
         SubCellInst_LFInst_8_LFInst_2_n1 ,
         SubCellInst_LFInst_8_LFInst_1_n7 ,
         SubCellInst_LFInst_8_LFInst_1_n6 ,
         SubCellInst_LFInst_8_LFInst_1_n5 ,
         SubCellInst_LFInst_8_LFInst_1_n4 ,
         SubCellInst_LFInst_8_LFInst_1_n3 ,
         SubCellInst_LFInst_8_LFInst_1_n2 ,
         SubCellInst_LFInst_8_LFInst_1_n1 ,
         SubCellInst_LFInst_8_LFInst_0_n2 ,
         SubCellInst_LFInst_8_LFInst_0_n1 ,
         SubCellInst_LFInst_9_LFInst_3_n8 ,
         SubCellInst_LFInst_9_LFInst_3_n7 ,
         SubCellInst_LFInst_9_LFInst_3_n6 ,
         SubCellInst_LFInst_9_LFInst_3_n5 ,
         SubCellInst_LFInst_9_LFInst_3_n4 ,
         SubCellInst_LFInst_9_LFInst_3_n3 ,
         SubCellInst_LFInst_9_LFInst_3_n2 ,
         SubCellInst_LFInst_9_LFInst_3_n1 ,
         SubCellInst_LFInst_9_LFInst_2_n10 ,
         SubCellInst_LFInst_9_LFInst_2_n9 ,
         SubCellInst_LFInst_9_LFInst_2_n8 ,
         SubCellInst_LFInst_9_LFInst_2_n7 ,
         SubCellInst_LFInst_9_LFInst_2_n6 ,
         SubCellInst_LFInst_9_LFInst_2_n5 ,
         SubCellInst_LFInst_9_LFInst_2_n4 ,
         SubCellInst_LFInst_9_LFInst_2_n3 ,
         SubCellInst_LFInst_9_LFInst_2_n2 ,
         SubCellInst_LFInst_9_LFInst_2_n1 ,
         SubCellInst_LFInst_9_LFInst_1_n7 ,
         SubCellInst_LFInst_9_LFInst_1_n6 ,
         SubCellInst_LFInst_9_LFInst_1_n5 ,
         SubCellInst_LFInst_9_LFInst_1_n4 ,
         SubCellInst_LFInst_9_LFInst_1_n3 ,
         SubCellInst_LFInst_9_LFInst_1_n2 ,
         SubCellInst_LFInst_9_LFInst_1_n1 ,
         SubCellInst_LFInst_9_LFInst_0_n2 ,
         SubCellInst_LFInst_9_LFInst_0_n1 ,
         SubCellInst_LFInst_10_LFInst_3_n8 ,
         SubCellInst_LFInst_10_LFInst_3_n7 ,
         SubCellInst_LFInst_10_LFInst_3_n6 ,
         SubCellInst_LFInst_10_LFInst_3_n5 ,
         SubCellInst_LFInst_10_LFInst_3_n4 ,
         SubCellInst_LFInst_10_LFInst_3_n3 ,
         SubCellInst_LFInst_10_LFInst_3_n2 ,
         SubCellInst_LFInst_10_LFInst_3_n1 ,
         SubCellInst_LFInst_10_LFInst_2_n10 ,
         SubCellInst_LFInst_10_LFInst_2_n9 ,
         SubCellInst_LFInst_10_LFInst_2_n8 ,
         SubCellInst_LFInst_10_LFInst_2_n7 ,
         SubCellInst_LFInst_10_LFInst_2_n6 ,
         SubCellInst_LFInst_10_LFInst_2_n5 ,
         SubCellInst_LFInst_10_LFInst_2_n4 ,
         SubCellInst_LFInst_10_LFInst_2_n3 ,
         SubCellInst_LFInst_10_LFInst_2_n2 ,
         SubCellInst_LFInst_10_LFInst_2_n1 ,
         SubCellInst_LFInst_10_LFInst_1_n7 ,
         SubCellInst_LFInst_10_LFInst_1_n6 ,
         SubCellInst_LFInst_10_LFInst_1_n5 ,
         SubCellInst_LFInst_10_LFInst_1_n4 ,
         SubCellInst_LFInst_10_LFInst_1_n3 ,
         SubCellInst_LFInst_10_LFInst_1_n2 ,
         SubCellInst_LFInst_10_LFInst_1_n1 ,
         SubCellInst_LFInst_10_LFInst_0_n2 ,
         SubCellInst_LFInst_10_LFInst_0_n1 ,
         SubCellInst_LFInst_11_LFInst_3_n8 ,
         SubCellInst_LFInst_11_LFInst_3_n7 ,
         SubCellInst_LFInst_11_LFInst_3_n6 ,
         SubCellInst_LFInst_11_LFInst_3_n5 ,
         SubCellInst_LFInst_11_LFInst_3_n4 ,
         SubCellInst_LFInst_11_LFInst_3_n3 ,
         SubCellInst_LFInst_11_LFInst_3_n2 ,
         SubCellInst_LFInst_11_LFInst_3_n1 ,
         SubCellInst_LFInst_11_LFInst_2_n10 ,
         SubCellInst_LFInst_11_LFInst_2_n9 ,
         SubCellInst_LFInst_11_LFInst_2_n8 ,
         SubCellInst_LFInst_11_LFInst_2_n7 ,
         SubCellInst_LFInst_11_LFInst_2_n6 ,
         SubCellInst_LFInst_11_LFInst_2_n5 ,
         SubCellInst_LFInst_11_LFInst_2_n4 ,
         SubCellInst_LFInst_11_LFInst_2_n3 ,
         SubCellInst_LFInst_11_LFInst_2_n2 ,
         SubCellInst_LFInst_11_LFInst_2_n1 ,
         SubCellInst_LFInst_11_LFInst_1_n7 ,
         SubCellInst_LFInst_11_LFInst_1_n6 ,
         SubCellInst_LFInst_11_LFInst_1_n5 ,
         SubCellInst_LFInst_11_LFInst_1_n4 ,
         SubCellInst_LFInst_11_LFInst_1_n3 ,
         SubCellInst_LFInst_11_LFInst_1_n2 ,
         SubCellInst_LFInst_11_LFInst_1_n1 ,
         SubCellInst_LFInst_11_LFInst_0_n2 ,
         SubCellInst_LFInst_11_LFInst_0_n1 ,
         SubCellInst_LFInst_12_LFInst_3_n8 ,
         SubCellInst_LFInst_12_LFInst_3_n7 ,
         SubCellInst_LFInst_12_LFInst_3_n6 ,
         SubCellInst_LFInst_12_LFInst_3_n5 ,
         SubCellInst_LFInst_12_LFInst_3_n4 ,
         SubCellInst_LFInst_12_LFInst_3_n3 ,
         SubCellInst_LFInst_12_LFInst_3_n2 ,
         SubCellInst_LFInst_12_LFInst_3_n1 ,
         SubCellInst_LFInst_12_LFInst_2_n10 ,
         SubCellInst_LFInst_12_LFInst_2_n9 ,
         SubCellInst_LFInst_12_LFInst_2_n8 ,
         SubCellInst_LFInst_12_LFInst_2_n7 ,
         SubCellInst_LFInst_12_LFInst_2_n6 ,
         SubCellInst_LFInst_12_LFInst_2_n5 ,
         SubCellInst_LFInst_12_LFInst_2_n4 ,
         SubCellInst_LFInst_12_LFInst_2_n3 ,
         SubCellInst_LFInst_12_LFInst_2_n2 ,
         SubCellInst_LFInst_12_LFInst_2_n1 ,
         SubCellInst_LFInst_12_LFInst_1_n7 ,
         SubCellInst_LFInst_12_LFInst_1_n6 ,
         SubCellInst_LFInst_12_LFInst_1_n5 ,
         SubCellInst_LFInst_12_LFInst_1_n4 ,
         SubCellInst_LFInst_12_LFInst_1_n3 ,
         SubCellInst_LFInst_12_LFInst_1_n2 ,
         SubCellInst_LFInst_12_LFInst_1_n1 ,
         SubCellInst_LFInst_12_LFInst_0_n2 ,
         SubCellInst_LFInst_12_LFInst_0_n1 ,
         SubCellInst_LFInst_13_LFInst_3_n8 ,
         SubCellInst_LFInst_13_LFInst_3_n7 ,
         SubCellInst_LFInst_13_LFInst_3_n6 ,
         SubCellInst_LFInst_13_LFInst_3_n5 ,
         SubCellInst_LFInst_13_LFInst_3_n4 ,
         SubCellInst_LFInst_13_LFInst_3_n3 ,
         SubCellInst_LFInst_13_LFInst_3_n2 ,
         SubCellInst_LFInst_13_LFInst_3_n1 ,
         SubCellInst_LFInst_13_LFInst_2_n10 ,
         SubCellInst_LFInst_13_LFInst_2_n9 ,
         SubCellInst_LFInst_13_LFInst_2_n8 ,
         SubCellInst_LFInst_13_LFInst_2_n7 ,
         SubCellInst_LFInst_13_LFInst_2_n6 ,
         SubCellInst_LFInst_13_LFInst_2_n5 ,
         SubCellInst_LFInst_13_LFInst_2_n4 ,
         SubCellInst_LFInst_13_LFInst_2_n3 ,
         SubCellInst_LFInst_13_LFInst_2_n2 ,
         SubCellInst_LFInst_13_LFInst_2_n1 ,
         SubCellInst_LFInst_13_LFInst_1_n7 ,
         SubCellInst_LFInst_13_LFInst_1_n6 ,
         SubCellInst_LFInst_13_LFInst_1_n5 ,
         SubCellInst_LFInst_13_LFInst_1_n4 ,
         SubCellInst_LFInst_13_LFInst_1_n3 ,
         SubCellInst_LFInst_13_LFInst_1_n2 ,
         SubCellInst_LFInst_13_LFInst_1_n1 ,
         SubCellInst_LFInst_13_LFInst_0_n2 ,
         SubCellInst_LFInst_13_LFInst_0_n1 ,
         SubCellInst_LFInst_14_LFInst_3_n8 ,
         SubCellInst_LFInst_14_LFInst_3_n7 ,
         SubCellInst_LFInst_14_LFInst_3_n6 ,
         SubCellInst_LFInst_14_LFInst_3_n5 ,
         SubCellInst_LFInst_14_LFInst_3_n4 ,
         SubCellInst_LFInst_14_LFInst_3_n3 ,
         SubCellInst_LFInst_14_LFInst_3_n2 ,
         SubCellInst_LFInst_14_LFInst_3_n1 ,
         SubCellInst_LFInst_14_LFInst_2_n10 ,
         SubCellInst_LFInst_14_LFInst_2_n9 ,
         SubCellInst_LFInst_14_LFInst_2_n8 ,
         SubCellInst_LFInst_14_LFInst_2_n7 ,
         SubCellInst_LFInst_14_LFInst_2_n6 ,
         SubCellInst_LFInst_14_LFInst_2_n5 ,
         SubCellInst_LFInst_14_LFInst_2_n4 ,
         SubCellInst_LFInst_14_LFInst_2_n3 ,
         SubCellInst_LFInst_14_LFInst_2_n2 ,
         SubCellInst_LFInst_14_LFInst_2_n1 ,
         SubCellInst_LFInst_14_LFInst_1_n7 ,
         SubCellInst_LFInst_14_LFInst_1_n6 ,
         SubCellInst_LFInst_14_LFInst_1_n5 ,
         SubCellInst_LFInst_14_LFInst_1_n4 ,
         SubCellInst_LFInst_14_LFInst_1_n3 ,
         SubCellInst_LFInst_14_LFInst_1_n2 ,
         SubCellInst_LFInst_14_LFInst_1_n1 ,
         SubCellInst_LFInst_14_LFInst_0_n2 ,
         SubCellInst_LFInst_14_LFInst_0_n1 ,
         SubCellInst_LFInst_15_LFInst_3_n8 ,
         SubCellInst_LFInst_15_LFInst_3_n7 ,
         SubCellInst_LFInst_15_LFInst_3_n6 ,
         SubCellInst_LFInst_15_LFInst_3_n5 ,
         SubCellInst_LFInst_15_LFInst_3_n4 ,
         SubCellInst_LFInst_15_LFInst_3_n3 ,
         SubCellInst_LFInst_15_LFInst_3_n2 ,
         SubCellInst_LFInst_15_LFInst_3_n1 ,
         SubCellInst_LFInst_15_LFInst_2_n10 ,
         SubCellInst_LFInst_15_LFInst_2_n9 ,
         SubCellInst_LFInst_15_LFInst_2_n8 ,
         SubCellInst_LFInst_15_LFInst_2_n7 ,
         SubCellInst_LFInst_15_LFInst_2_n6 ,
         SubCellInst_LFInst_15_LFInst_2_n5 ,
         SubCellInst_LFInst_15_LFInst_2_n4 ,
         SubCellInst_LFInst_15_LFInst_2_n3 ,
         SubCellInst_LFInst_15_LFInst_2_n2 ,
         SubCellInst_LFInst_15_LFInst_2_n1 ,
         SubCellInst_LFInst_15_LFInst_1_n7 ,
         SubCellInst_LFInst_15_LFInst_1_n6 ,
         SubCellInst_LFInst_15_LFInst_1_n5 ,
         SubCellInst_LFInst_15_LFInst_1_n4 ,
         SubCellInst_LFInst_15_LFInst_1_n3 ,
         SubCellInst_LFInst_15_LFInst_1_n2 ,
         SubCellInst_LFInst_15_LFInst_1_n1 ,
         SubCellInst_LFInst_15_LFInst_0_n2 ,
         SubCellInst_LFInst_15_LFInst_0_n1 , MCInst1_MC0_v0_2Inst_0_n1 ,
         MCInst1_MC0_v1_2Inst_0_n1 , MCInst1_MC0_v2_3Inst_0_n2 ,
         MCInst1_MC0_v2_3Inst_0_n1 , MCInst1_MC0_v3_3Inst_0_n1 ,
         MCInst1_MC0_v0_2Inst_1_n1 , MCInst1_MC0_v2_1Inst_1_n1 ,
         MCInst1_MC0_v2_2Inst_1_n2 , MCInst1_MC0_v2_2Inst_1_n1 ,
         MCInst1_MC0_v3_3Inst_1_n1 , MCInst1_MC0_v1_1Inst_2_n1 ,
         MCInst1_MC0_v1_2Inst_2_n1 , MCInst1_MC0_v2_1Inst_2_n1 ,
         MCInst1_MC0_v2_2Inst_2_n1 , MCInst1_MC0_v3_1Inst_2_n1 ,
         MCInst1_MC0_v1_2Inst_3_n2 , MCInst1_MC0_v1_2Inst_3_n1 ,
         MCInst1_MC0_v2_2Inst_3_n1 , MCInst1_MC0_v2_3Inst_3_n1 ,
         MCInst1_MC0_r0Inst_XORInst_0_0_n3 ,
         MCInst1_MC0_r0Inst_XORInst_0_0_n2 ,
         MCInst1_MC0_r0Inst_XORInst_0_0_n1 ,
         MCInst1_MC0_r0Inst_XORInst_0_1_n6 ,
         MCInst1_MC0_r0Inst_XORInst_0_1_n5 ,
         MCInst1_MC0_r0Inst_XORInst_0_1_n4 ,
         MCInst1_MC0_r0Inst_XORInst_0_2_n6 ,
         MCInst1_MC0_r0Inst_XORInst_0_2_n5 ,
         MCInst1_MC0_r0Inst_XORInst_0_2_n4 ,
         MCInst1_MC0_r0Inst_XORInst_0_3_n6 ,
         MCInst1_MC0_r0Inst_XORInst_0_3_n5 ,
         MCInst1_MC0_r0Inst_XORInst_0_3_n4 ,
         MCInst1_MC0_r1Inst_XORInst_0_0_n6 ,
         MCInst1_MC0_r1Inst_XORInst_0_0_n5 ,
         MCInst1_MC0_r1Inst_XORInst_0_0_n4 ,
         MCInst1_MC0_r1Inst_XORInst_0_1_n6 ,
         MCInst1_MC0_r1Inst_XORInst_0_1_n5 ,
         MCInst1_MC0_r1Inst_XORInst_0_1_n4 ,
         MCInst1_MC0_r1Inst_XORInst_0_2_n6 ,
         MCInst1_MC0_r1Inst_XORInst_0_2_n5 ,
         MCInst1_MC0_r1Inst_XORInst_0_2_n4 ,
         MCInst1_MC0_r1Inst_XORInst_0_3_n6 ,
         MCInst1_MC0_r1Inst_XORInst_0_3_n5 ,
         MCInst1_MC0_r1Inst_XORInst_0_3_n4 ,
         MCInst1_MC0_r2Inst_XORInst_0_0_n6 ,
         MCInst1_MC0_r2Inst_XORInst_0_0_n5 ,
         MCInst1_MC0_r2Inst_XORInst_0_0_n4 ,
         MCInst1_MC0_r2Inst_XORInst_0_1_n6 ,
         MCInst1_MC0_r2Inst_XORInst_0_1_n5 ,
         MCInst1_MC0_r2Inst_XORInst_0_1_n4 ,
         MCInst1_MC0_r2Inst_XORInst_0_2_n6 ,
         MCInst1_MC0_r2Inst_XORInst_0_2_n5 ,
         MCInst1_MC0_r2Inst_XORInst_0_2_n4 ,
         MCInst1_MC0_r2Inst_XORInst_0_3_n6 ,
         MCInst1_MC0_r2Inst_XORInst_0_3_n5 ,
         MCInst1_MC0_r2Inst_XORInst_0_3_n4 ,
         MCInst1_MC0_r3Inst_XORInst_0_0_n6 ,
         MCInst1_MC0_r3Inst_XORInst_0_0_n5 ,
         MCInst1_MC0_r3Inst_XORInst_0_0_n4 ,
         MCInst1_MC0_r3Inst_XORInst_0_1_n6 ,
         MCInst1_MC0_r3Inst_XORInst_0_1_n5 ,
         MCInst1_MC0_r3Inst_XORInst_0_1_n4 ,
         MCInst1_MC0_r3Inst_XORInst_0_2_n6 ,
         MCInst1_MC0_r3Inst_XORInst_0_2_n5 ,
         MCInst1_MC0_r3Inst_XORInst_0_2_n4 ,
         MCInst1_MC0_r3Inst_XORInst_0_3_n6 ,
         MCInst1_MC0_r3Inst_XORInst_0_3_n5 ,
         MCInst1_MC0_r3Inst_XORInst_0_3_n4 , MCInst1_MC1_v0_2Inst_0_n1 ,
         MCInst1_MC1_v1_2Inst_0_n1 , MCInst1_MC1_v2_3Inst_0_n2 ,
         MCInst1_MC1_v2_3Inst_0_n1 , MCInst1_MC1_v3_3Inst_0_n1 ,
         MCInst1_MC1_v0_2Inst_1_n1 , MCInst1_MC1_v2_1Inst_1_n1 ,
         MCInst1_MC1_v2_2Inst_1_n2 , MCInst1_MC1_v2_2Inst_1_n1 ,
         MCInst1_MC1_v3_3Inst_1_n1 , MCInst1_MC1_v1_1Inst_2_n1 ,
         MCInst1_MC1_v1_2Inst_2_n1 , MCInst1_MC1_v2_1Inst_2_n1 ,
         MCInst1_MC1_v2_2Inst_2_n1 , MCInst1_MC1_v3_1Inst_2_n1 ,
         MCInst1_MC1_v1_2Inst_3_n2 , MCInst1_MC1_v1_2Inst_3_n1 ,
         MCInst1_MC1_v2_2Inst_3_n1 , MCInst1_MC1_v2_3Inst_3_n1 ,
         MCInst1_MC1_r0Inst_XORInst_0_0_n6 ,
         MCInst1_MC1_r0Inst_XORInst_0_0_n5 ,
         MCInst1_MC1_r0Inst_XORInst_0_0_n4 ,
         MCInst1_MC1_r0Inst_XORInst_0_1_n6 ,
         MCInst1_MC1_r0Inst_XORInst_0_1_n5 ,
         MCInst1_MC1_r0Inst_XORInst_0_1_n4 ,
         MCInst1_MC1_r0Inst_XORInst_0_2_n6 ,
         MCInst1_MC1_r0Inst_XORInst_0_2_n5 ,
         MCInst1_MC1_r0Inst_XORInst_0_2_n4 ,
         MCInst1_MC1_r0Inst_XORInst_0_3_n6 ,
         MCInst1_MC1_r0Inst_XORInst_0_3_n5 ,
         MCInst1_MC1_r0Inst_XORInst_0_3_n4 ,
         MCInst1_MC1_r1Inst_XORInst_0_0_n6 ,
         MCInst1_MC1_r1Inst_XORInst_0_0_n5 ,
         MCInst1_MC1_r1Inst_XORInst_0_0_n4 ,
         MCInst1_MC1_r1Inst_XORInst_0_1_n6 ,
         MCInst1_MC1_r1Inst_XORInst_0_1_n5 ,
         MCInst1_MC1_r1Inst_XORInst_0_1_n4 ,
         MCInst1_MC1_r1Inst_XORInst_0_2_n6 ,
         MCInst1_MC1_r1Inst_XORInst_0_2_n5 ,
         MCInst1_MC1_r1Inst_XORInst_0_2_n4 ,
         MCInst1_MC1_r1Inst_XORInst_0_3_n6 ,
         MCInst1_MC1_r1Inst_XORInst_0_3_n5 ,
         MCInst1_MC1_r1Inst_XORInst_0_3_n4 ,
         MCInst1_MC1_r2Inst_XORInst_0_0_n6 ,
         MCInst1_MC1_r2Inst_XORInst_0_0_n5 ,
         MCInst1_MC1_r2Inst_XORInst_0_0_n4 ,
         MCInst1_MC1_r2Inst_XORInst_0_1_n6 ,
         MCInst1_MC1_r2Inst_XORInst_0_1_n5 ,
         MCInst1_MC1_r2Inst_XORInst_0_1_n4 ,
         MCInst1_MC1_r2Inst_XORInst_0_2_n6 ,
         MCInst1_MC1_r2Inst_XORInst_0_2_n5 ,
         MCInst1_MC1_r2Inst_XORInst_0_2_n4 ,
         MCInst1_MC1_r2Inst_XORInst_0_3_n6 ,
         MCInst1_MC1_r2Inst_XORInst_0_3_n5 ,
         MCInst1_MC1_r2Inst_XORInst_0_3_n4 ,
         MCInst1_MC1_r3Inst_XORInst_0_0_n6 ,
         MCInst1_MC1_r3Inst_XORInst_0_0_n5 ,
         MCInst1_MC1_r3Inst_XORInst_0_0_n4 ,
         MCInst1_MC1_r3Inst_XORInst_0_1_n6 ,
         MCInst1_MC1_r3Inst_XORInst_0_1_n5 ,
         MCInst1_MC1_r3Inst_XORInst_0_1_n4 ,
         MCInst1_MC1_r3Inst_XORInst_0_2_n6 ,
         MCInst1_MC1_r3Inst_XORInst_0_2_n5 ,
         MCInst1_MC1_r3Inst_XORInst_0_2_n4 ,
         MCInst1_MC1_r3Inst_XORInst_0_3_n6 ,
         MCInst1_MC1_r3Inst_XORInst_0_3_n5 ,
         MCInst1_MC1_r3Inst_XORInst_0_3_n4 , MCInst1_MC2_v0_2Inst_0_n1 ,
         MCInst1_MC2_v1_2Inst_0_n1 , MCInst1_MC2_v2_3Inst_0_n2 ,
         MCInst1_MC2_v2_3Inst_0_n1 , MCInst1_MC2_v3_3Inst_0_n1 ,
         MCInst1_MC2_v0_2Inst_1_n1 , MCInst1_MC2_v2_1Inst_1_n1 ,
         MCInst1_MC2_v2_2Inst_1_n2 , MCInst1_MC2_v2_2Inst_1_n1 ,
         MCInst1_MC2_v3_3Inst_1_n1 , MCInst1_MC2_v1_1Inst_2_n1 ,
         MCInst1_MC2_v1_2Inst_2_n1 , MCInst1_MC2_v2_1Inst_2_n1 ,
         MCInst1_MC2_v2_2Inst_2_n1 , MCInst1_MC2_v3_1Inst_2_n1 ,
         MCInst1_MC2_v1_2Inst_3_n2 , MCInst1_MC2_v1_2Inst_3_n1 ,
         MCInst1_MC2_v2_2Inst_3_n1 , MCInst1_MC2_v2_3Inst_3_n1 ,
         MCInst1_MC2_r0Inst_XORInst_0_0_n6 ,
         MCInst1_MC2_r0Inst_XORInst_0_0_n5 ,
         MCInst1_MC2_r0Inst_XORInst_0_0_n4 ,
         MCInst1_MC2_r0Inst_XORInst_0_1_n6 ,
         MCInst1_MC2_r0Inst_XORInst_0_1_n5 ,
         MCInst1_MC2_r0Inst_XORInst_0_1_n4 ,
         MCInst1_MC2_r0Inst_XORInst_0_2_n6 ,
         MCInst1_MC2_r0Inst_XORInst_0_2_n5 ,
         MCInst1_MC2_r0Inst_XORInst_0_2_n4 ,
         MCInst1_MC2_r0Inst_XORInst_0_3_n6 ,
         MCInst1_MC2_r0Inst_XORInst_0_3_n5 ,
         MCInst1_MC2_r0Inst_XORInst_0_3_n4 ,
         MCInst1_MC2_r1Inst_XORInst_0_0_n6 ,
         MCInst1_MC2_r1Inst_XORInst_0_0_n5 ,
         MCInst1_MC2_r1Inst_XORInst_0_0_n4 ,
         MCInst1_MC2_r1Inst_XORInst_0_1_n6 ,
         MCInst1_MC2_r1Inst_XORInst_0_1_n5 ,
         MCInst1_MC2_r1Inst_XORInst_0_1_n4 ,
         MCInst1_MC2_r1Inst_XORInst_0_2_n6 ,
         MCInst1_MC2_r1Inst_XORInst_0_2_n5 ,
         MCInst1_MC2_r1Inst_XORInst_0_2_n4 ,
         MCInst1_MC2_r1Inst_XORInst_0_3_n6 ,
         MCInst1_MC2_r1Inst_XORInst_0_3_n5 ,
         MCInst1_MC2_r1Inst_XORInst_0_3_n4 ,
         MCInst1_MC2_r2Inst_XORInst_0_0_n6 ,
         MCInst1_MC2_r2Inst_XORInst_0_0_n5 ,
         MCInst1_MC2_r2Inst_XORInst_0_0_n4 ,
         MCInst1_MC2_r2Inst_XORInst_0_1_n6 ,
         MCInst1_MC2_r2Inst_XORInst_0_1_n5 ,
         MCInst1_MC2_r2Inst_XORInst_0_1_n4 ,
         MCInst1_MC2_r2Inst_XORInst_0_2_n6 ,
         MCInst1_MC2_r2Inst_XORInst_0_2_n5 ,
         MCInst1_MC2_r2Inst_XORInst_0_2_n4 ,
         MCInst1_MC2_r2Inst_XORInst_0_3_n6 ,
         MCInst1_MC2_r2Inst_XORInst_0_3_n5 ,
         MCInst1_MC2_r2Inst_XORInst_0_3_n4 ,
         MCInst1_MC2_r3Inst_XORInst_0_0_n6 ,
         MCInst1_MC2_r3Inst_XORInst_0_0_n5 ,
         MCInst1_MC2_r3Inst_XORInst_0_0_n4 ,
         MCInst1_MC2_r3Inst_XORInst_0_1_n6 ,
         MCInst1_MC2_r3Inst_XORInst_0_1_n5 ,
         MCInst1_MC2_r3Inst_XORInst_0_1_n4 ,
         MCInst1_MC2_r3Inst_XORInst_0_2_n6 ,
         MCInst1_MC2_r3Inst_XORInst_0_2_n5 ,
         MCInst1_MC2_r3Inst_XORInst_0_2_n4 ,
         MCInst1_MC2_r3Inst_XORInst_0_3_n6 ,
         MCInst1_MC2_r3Inst_XORInst_0_3_n5 ,
         MCInst1_MC2_r3Inst_XORInst_0_3_n4 , MCInst1_MC3_v0_2Inst_0_n1 ,
         MCInst1_MC3_v1_2Inst_0_n1 , MCInst1_MC3_v2_3Inst_0_n2 ,
         MCInst1_MC3_v2_3Inst_0_n1 , MCInst1_MC3_v3_3Inst_0_n1 ,
         MCInst1_MC3_v0_2Inst_1_n1 , MCInst1_MC3_v2_1Inst_1_n1 ,
         MCInst1_MC3_v2_2Inst_1_n2 , MCInst1_MC3_v2_2Inst_1_n1 ,
         MCInst1_MC3_v3_3Inst_1_n1 , MCInst1_MC3_v1_1Inst_2_n1 ,
         MCInst1_MC3_v1_2Inst_2_n1 , MCInst1_MC3_v2_1Inst_2_n1 ,
         MCInst1_MC3_v2_2Inst_2_n1 , MCInst1_MC3_v3_1Inst_2_n1 ,
         MCInst1_MC3_v1_2Inst_3_n2 , MCInst1_MC3_v1_2Inst_3_n1 ,
         MCInst1_MC3_v2_2Inst_3_n1 , MCInst1_MC3_v2_3Inst_3_n1 ,
         MCInst1_MC3_r0Inst_XORInst_0_0_n6 ,
         MCInst1_MC3_r0Inst_XORInst_0_0_n5 ,
         MCInst1_MC3_r0Inst_XORInst_0_0_n4 ,
         MCInst1_MC3_r0Inst_XORInst_0_1_n6 ,
         MCInst1_MC3_r0Inst_XORInst_0_1_n5 ,
         MCInst1_MC3_r0Inst_XORInst_0_1_n4 ,
         MCInst1_MC3_r0Inst_XORInst_0_2_n6 ,
         MCInst1_MC3_r0Inst_XORInst_0_2_n5 ,
         MCInst1_MC3_r0Inst_XORInst_0_2_n4 ,
         MCInst1_MC3_r0Inst_XORInst_0_3_n6 ,
         MCInst1_MC3_r0Inst_XORInst_0_3_n5 ,
         MCInst1_MC3_r0Inst_XORInst_0_3_n4 ,
         MCInst1_MC3_r1Inst_XORInst_0_0_n6 ,
         MCInst1_MC3_r1Inst_XORInst_0_0_n5 ,
         MCInst1_MC3_r1Inst_XORInst_0_0_n4 ,
         MCInst1_MC3_r1Inst_XORInst_0_1_n6 ,
         MCInst1_MC3_r1Inst_XORInst_0_1_n5 ,
         MCInst1_MC3_r1Inst_XORInst_0_1_n4 ,
         MCInst1_MC3_r1Inst_XORInst_0_2_n6 ,
         MCInst1_MC3_r1Inst_XORInst_0_2_n5 ,
         MCInst1_MC3_r1Inst_XORInst_0_2_n4 ,
         MCInst1_MC3_r1Inst_XORInst_0_3_n6 ,
         MCInst1_MC3_r1Inst_XORInst_0_3_n5 ,
         MCInst1_MC3_r1Inst_XORInst_0_3_n4 ,
         MCInst1_MC3_r2Inst_XORInst_0_0_n6 ,
         MCInst1_MC3_r2Inst_XORInst_0_0_n5 ,
         MCInst1_MC3_r2Inst_XORInst_0_0_n4 ,
         MCInst1_MC3_r2Inst_XORInst_0_1_n6 ,
         MCInst1_MC3_r2Inst_XORInst_0_1_n5 ,
         MCInst1_MC3_r2Inst_XORInst_0_1_n4 ,
         MCInst1_MC3_r2Inst_XORInst_0_2_n6 ,
         MCInst1_MC3_r2Inst_XORInst_0_2_n5 ,
         MCInst1_MC3_r2Inst_XORInst_0_2_n4 ,
         MCInst1_MC3_r2Inst_XORInst_0_3_n6 ,
         MCInst1_MC3_r2Inst_XORInst_0_3_n5 ,
         MCInst1_MC3_r2Inst_XORInst_0_3_n4 ,
         MCInst1_MC3_r3Inst_XORInst_0_0_n6 ,
         MCInst1_MC3_r3Inst_XORInst_0_0_n5 ,
         MCInst1_MC3_r3Inst_XORInst_0_0_n4 ,
         MCInst1_MC3_r3Inst_XORInst_0_1_n6 ,
         MCInst1_MC3_r3Inst_XORInst_0_1_n5 ,
         MCInst1_MC3_r3Inst_XORInst_0_1_n4 ,
         MCInst1_MC3_r3Inst_XORInst_0_2_n6 ,
         MCInst1_MC3_r3Inst_XORInst_0_2_n5 ,
         MCInst1_MC3_r3Inst_XORInst_0_2_n4 ,
         MCInst1_MC3_r3Inst_XORInst_0_3_n6 ,
         MCInst1_MC3_r3Inst_XORInst_0_3_n5 ,
         MCInst1_MC3_r3Inst_XORInst_0_3_n4 , FSMMUX_MUXInst_0_n2 ,
         FSMMUX_MUXInst_0_n1 , FSMMUX_MUXInst_1_n2 , FSMMUX_MUXInst_1_n1 ,
         FSMMUX_MUXInst_2_n2 , FSMMUX_MUXInst_2_n1 , FSMMUX_MUXInst_3_n2 ,
         FSMMUX_MUXInst_3_n1 , FSMMUX_MUXInst_4_n2 , FSMMUX_MUXInst_4_n1 ,
         FSMMUX_MUXInst_5_n2 , FSMMUX_MUXInst_5_n1 ,
         FSMUpdateInst_StateUpdateInst_0_n6 ,
         FSMUpdateInst_StateUpdateInst_0_n5 ,
         FSMUpdateInst_StateUpdateInst_0_n4 ,
         FSMUpdateInst_StateUpdateInst_0_n3 ,
         FSMUpdateInst_StateUpdateInst_0_n2 ,
         FSMUpdateInst_StateUpdateInst_0_n1 ,
         FSMUpdateInst_StateUpdateInst_2_n4 ,
         FSMUpdateInst_StateUpdateInst_2_n3 ,
         FSMUpdateInst_StateUpdateInst_2_n2 ,
         FSMUpdateInst_StateUpdateInst_2_n1 ,
         FSMUpdateInst_StateUpdateInst_5_n4 ,
         FSMUpdateInst_StateUpdateInst_5_n3 ,
         FSMUpdateInst_StateUpdateInst_5_n2 ,
         FSMUpdateInst_StateUpdateInst_5_n1 , FSMSignalsInst_AddKeyInst_n14 ,
         FSMSignalsInst_AddKeyInst_n13 , FSMSignalsInst_AddKeyInst_n12 ,
         FSMSignalsInst_AddKeyInst_n11 , FSMSignalsInst_AddKeyInst_n10 ,
         FSMSignalsInst_AddKeyInst_n9 , FSMSignalsInst_AddKeyInst_n8 ,
         FSMSignalsInst_AddKeyInst_n7 , FSMSignalsInst_AddKeyInst_n6 ,
         FSMSignalsInst_AddKeyInst_n5 , FSMSignalsInst_AddKeyInst_n4 ,
         FSMSignalsInst_AddKeyInst_n3 , FSMSignalsInst_AddKeyInst_n2 ,
         FSMSignalsInst_AddKeyInst_n1 , FSMSignalsInst_doneInst_n4 ,
         FSMSignalsInst_doneInst_n3 , FSMSignalsInst_doneInst_n2 ,
         FSMSignalsInst_doneInst_n1 ;
  wire   [63:0] Feedback;
  wire   [63:0] StateRegInput;
  wire   [63:0] StateRegOutput;
  wire   [63:0] AddKeyMUXOutput;
  wire   [5:0] FSM;
  wire   [31:0] AddConstOutput;
  wire   [63:0] ShiftRowsOutput;
  wire   [5:0] FSMUpdate;
  wire   [5:0] FSMSelected;
  wire   [3:0] MCInst1_MC0_v3_3 ;
  wire   [3:0] MCInst1_MC0_v3_2 ;
  wire   [3:0] MCInst1_MC0_v3_1 ;
  wire   [3:0] MCInst1_MC0_v3_0 ;
  wire   [3:0] MCInst1_MC0_v2_3 ;
  wire   [3:0] MCInst1_MC0_v2_2 ;
  wire   [3:0] MCInst1_MC0_v2_1 ;
  wire   [3:0] MCInst1_MC0_v2_0 ;
  wire   [3:0] MCInst1_MC0_v1_3 ;
  wire   [3:0] MCInst1_MC0_v1_2 ;
  wire   [3:0] MCInst1_MC0_v1_1 ;
  wire   [3:0] MCInst1_MC0_v0_3 ;
  wire   [3:0] MCInst1_MC0_v0_2 ;
  wire   [3:0] MCInst1_MC0_v0_1 ;
  wire   [3:0] MCInst1_MC0_v0_0 ;
  wire   [3:0] MCInst1_MC1_v3_3 ;
  wire   [3:0] MCInst1_MC1_v3_2 ;
  wire   [3:0] MCInst1_MC1_v3_1 ;
  wire   [3:0] MCInst1_MC1_v3_0 ;
  wire   [3:0] MCInst1_MC1_v2_3 ;
  wire   [3:0] MCInst1_MC1_v2_2 ;
  wire   [3:0] MCInst1_MC1_v2_1 ;
  wire   [3:0] MCInst1_MC1_v2_0 ;
  wire   [3:0] MCInst1_MC1_v1_3 ;
  wire   [3:0] MCInst1_MC1_v1_2 ;
  wire   [3:0] MCInst1_MC1_v1_1 ;
  wire   [3:0] MCInst1_MC1_v0_3 ;
  wire   [3:0] MCInst1_MC1_v0_2 ;
  wire   [3:0] MCInst1_MC1_v0_1 ;
  wire   [3:0] MCInst1_MC1_v0_0 ;
  wire   [3:0] MCInst1_MC2_v3_3 ;
  wire   [3:0] MCInst1_MC2_v3_2 ;
  wire   [3:0] MCInst1_MC2_v3_1 ;
  wire   [3:0] MCInst1_MC2_v3_0 ;
  wire   [3:0] MCInst1_MC2_v2_3 ;
  wire   [3:0] MCInst1_MC2_v2_2 ;
  wire   [3:0] MCInst1_MC2_v2_1 ;
  wire   [3:0] MCInst1_MC2_v2_0 ;
  wire   [3:0] MCInst1_MC2_v1_3 ;
  wire   [3:0] MCInst1_MC2_v1_2 ;
  wire   [3:0] MCInst1_MC2_v1_1 ;
  wire   [3:0] MCInst1_MC2_v0_3 ;
  wire   [3:0] MCInst1_MC2_v0_2 ;
  wire   [3:0] MCInst1_MC2_v0_1 ;
  wire   [3:0] MCInst1_MC2_v0_0 ;
  wire   [3:0] MCInst1_MC3_v3_3 ;
  wire   [3:0] MCInst1_MC3_v3_2 ;
  wire   [3:0] MCInst1_MC3_v3_1 ;
  wire   [3:0] MCInst1_MC3_v3_0 ;
  wire   [3:0] MCInst1_MC3_v2_3 ;
  wire   [3:0] MCInst1_MC3_v2_2 ;
  wire   [3:0] MCInst1_MC3_v2_1 ;
  wire   [3:0] MCInst1_MC3_v2_0 ;
  wire   [3:0] MCInst1_MC3_v1_3 ;
  wire   [3:0] MCInst1_MC3_v1_2 ;
  wire   [3:0] MCInst1_MC3_v1_1 ;
  wire   [3:0] MCInst1_MC3_v0_3 ;
  wire   [3:0] MCInst1_MC3_v0_2 ;
  wire   [3:0] MCInst1_MC3_v0_1 ;
  wire   [3:0] MCInst1_MC3_v0_0 ;

  AND2 PlaintextMUX_MUXInst_0_U3  ( .A(Plaintext[0]), .B(rst), .Z(
        PlaintextMUX_MUXInst_0_n1 ) );
  ORN2 PlaintextMUX_MUXInst_0_U2  ( .A(rst), .B(Feedback[0]), .Z(
        PlaintextMUX_MUXInst_0_n2 ) );
  ORN2 PlaintextMUX_MUXInst_0_U1  ( .A(PlaintextMUX_MUXInst_0_n1 ), .B(
        PlaintextMUX_MUXInst_0_n2 ), .Z(StateRegInput[0]) );
  AND2 PlaintextMUX_MUXInst_1_U3  ( .A(Plaintext[1]), .B(rst), .Z(
        PlaintextMUX_MUXInst_1_n1 ) );
  ORN2 PlaintextMUX_MUXInst_1_U2  ( .A(rst), .B(Feedback[1]), .Z(
        PlaintextMUX_MUXInst_1_n2 ) );
  ORN2 PlaintextMUX_MUXInst_1_U1  ( .A(PlaintextMUX_MUXInst_1_n1 ), .B(
        PlaintextMUX_MUXInst_1_n2 ), .Z(StateRegInput[1]) );
  AND2 PlaintextMUX_MUXInst_2_U3  ( .A(Plaintext[2]), .B(rst), .Z(
        PlaintextMUX_MUXInst_2_n1 ) );
  ORN2 PlaintextMUX_MUXInst_2_U2  ( .A(rst), .B(Feedback[2]), .Z(
        PlaintextMUX_MUXInst_2_n2 ) );
  ORN2 PlaintextMUX_MUXInst_2_U1  ( .A(PlaintextMUX_MUXInst_2_n1 ), .B(
        PlaintextMUX_MUXInst_2_n2 ), .Z(StateRegInput[2]) );
  AND2 PlaintextMUX_MUXInst_3_U3  ( .A(Plaintext[3]), .B(rst), .Z(
        PlaintextMUX_MUXInst_3_n1 ) );
  ORN2 PlaintextMUX_MUXInst_3_U2  ( .A(rst), .B(Feedback[3]), .Z(
        PlaintextMUX_MUXInst_3_n2 ) );
  ORN2 PlaintextMUX_MUXInst_3_U1  ( .A(PlaintextMUX_MUXInst_3_n1 ), .B(
        PlaintextMUX_MUXInst_3_n2 ), .Z(StateRegInput[3]) );
  AND2 PlaintextMUX_MUXInst_4_U3  ( .A(Plaintext[4]), .B(rst), .Z(
        PlaintextMUX_MUXInst_4_n1 ) );
  ORN2 PlaintextMUX_MUXInst_4_U2  ( .A(rst), .B(Feedback[4]), .Z(
        PlaintextMUX_MUXInst_4_n2 ) );
  ORN2 PlaintextMUX_MUXInst_4_U1  ( .A(PlaintextMUX_MUXInst_4_n1 ), .B(
        PlaintextMUX_MUXInst_4_n2 ), .Z(StateRegInput[4]) );
  AND2 PlaintextMUX_MUXInst_5_U3  ( .A(Plaintext[5]), .B(rst), .Z(
        PlaintextMUX_MUXInst_5_n1 ) );
  ORN2 PlaintextMUX_MUXInst_5_U2  ( .A(rst), .B(Feedback[5]), .Z(
        PlaintextMUX_MUXInst_5_n2 ) );
  ORN2 PlaintextMUX_MUXInst_5_U1  ( .A(PlaintextMUX_MUXInst_5_n1 ), .B(
        PlaintextMUX_MUXInst_5_n2 ), .Z(StateRegInput[5]) );
  AND2 PlaintextMUX_MUXInst_6_U3  ( .A(Plaintext[6]), .B(rst), .Z(
        PlaintextMUX_MUXInst_6_n1 ) );
  ORN2 PlaintextMUX_MUXInst_6_U2  ( .A(rst), .B(Feedback[6]), .Z(
        PlaintextMUX_MUXInst_6_n2 ) );
  ORN2 PlaintextMUX_MUXInst_6_U1  ( .A(PlaintextMUX_MUXInst_6_n1 ), .B(
        PlaintextMUX_MUXInst_6_n2 ), .Z(StateRegInput[6]) );
  AND2 PlaintextMUX_MUXInst_7_U3  ( .A(Plaintext[7]), .B(rst), .Z(
        PlaintextMUX_MUXInst_7_n1 ) );
  ORN2 PlaintextMUX_MUXInst_7_U2  ( .A(rst), .B(Feedback[7]), .Z(
        PlaintextMUX_MUXInst_7_n2 ) );
  ORN2 PlaintextMUX_MUXInst_7_U1  ( .A(PlaintextMUX_MUXInst_7_n1 ), .B(
        PlaintextMUX_MUXInst_7_n2 ), .Z(StateRegInput[7]) );
  AND2 PlaintextMUX_MUXInst_8_U3  ( .A(Plaintext[8]), .B(rst), .Z(
        PlaintextMUX_MUXInst_8_n1 ) );
  ORN2 PlaintextMUX_MUXInst_8_U2  ( .A(rst), .B(Feedback[8]), .Z(
        PlaintextMUX_MUXInst_8_n2 ) );
  ORN2 PlaintextMUX_MUXInst_8_U1  ( .A(PlaintextMUX_MUXInst_8_n1 ), .B(
        PlaintextMUX_MUXInst_8_n2 ), .Z(StateRegInput[8]) );
  AND2 PlaintextMUX_MUXInst_9_U3  ( .A(Plaintext[9]), .B(rst), .Z(
        PlaintextMUX_MUXInst_9_n1 ) );
  ORN2 PlaintextMUX_MUXInst_9_U2  ( .A(rst), .B(Feedback[9]), .Z(
        PlaintextMUX_MUXInst_9_n2 ) );
  ORN2 PlaintextMUX_MUXInst_9_U1  ( .A(PlaintextMUX_MUXInst_9_n1 ), .B(
        PlaintextMUX_MUXInst_9_n2 ), .Z(StateRegInput[9]) );
  AND2 PlaintextMUX_MUXInst_10_U3  ( .A(Plaintext[10]), .B(rst), .Z(
        PlaintextMUX_MUXInst_10_n1 ) );
  ORN2 PlaintextMUX_MUXInst_10_U2  ( .A(rst), .B(Feedback[10]), .Z(
        PlaintextMUX_MUXInst_10_n2 ) );
  ORN2 PlaintextMUX_MUXInst_10_U1  ( .A(PlaintextMUX_MUXInst_10_n1 ), .B(
        PlaintextMUX_MUXInst_10_n2 ), .Z(StateRegInput[10]) );
  AND2 PlaintextMUX_MUXInst_11_U3  ( .A(Plaintext[11]), .B(rst), .Z(
        PlaintextMUX_MUXInst_11_n1 ) );
  ORN2 PlaintextMUX_MUXInst_11_U2  ( .A(rst), .B(Feedback[11]), .Z(
        PlaintextMUX_MUXInst_11_n2 ) );
  ORN2 PlaintextMUX_MUXInst_11_U1  ( .A(PlaintextMUX_MUXInst_11_n1 ), .B(
        PlaintextMUX_MUXInst_11_n2 ), .Z(StateRegInput[11]) );
  AND2 PlaintextMUX_MUXInst_12_U3  ( .A(Plaintext[12]), .B(rst), .Z(
        PlaintextMUX_MUXInst_12_n1 ) );
  ORN2 PlaintextMUX_MUXInst_12_U2  ( .A(rst), .B(Feedback[12]), .Z(
        PlaintextMUX_MUXInst_12_n2 ) );
  ORN2 PlaintextMUX_MUXInst_12_U1  ( .A(PlaintextMUX_MUXInst_12_n1 ), .B(
        PlaintextMUX_MUXInst_12_n2 ), .Z(StateRegInput[12]) );
  AND2 PlaintextMUX_MUXInst_13_U3  ( .A(Plaintext[13]), .B(rst), .Z(
        PlaintextMUX_MUXInst_13_n1 ) );
  ORN2 PlaintextMUX_MUXInst_13_U2  ( .A(rst), .B(Feedback[13]), .Z(
        PlaintextMUX_MUXInst_13_n2 ) );
  ORN2 PlaintextMUX_MUXInst_13_U1  ( .A(PlaintextMUX_MUXInst_13_n1 ), .B(
        PlaintextMUX_MUXInst_13_n2 ), .Z(StateRegInput[13]) );
  AND2 PlaintextMUX_MUXInst_14_U3  ( .A(Plaintext[14]), .B(rst), .Z(
        PlaintextMUX_MUXInst_14_n1 ) );
  ORN2 PlaintextMUX_MUXInst_14_U2  ( .A(rst), .B(Feedback[14]), .Z(
        PlaintextMUX_MUXInst_14_n2 ) );
  ORN2 PlaintextMUX_MUXInst_14_U1  ( .A(PlaintextMUX_MUXInst_14_n1 ), .B(
        PlaintextMUX_MUXInst_14_n2 ), .Z(StateRegInput[14]) );
  AND2 PlaintextMUX_MUXInst_15_U3  ( .A(Plaintext[15]), .B(rst), .Z(
        PlaintextMUX_MUXInst_15_n1 ) );
  ORN2 PlaintextMUX_MUXInst_15_U2  ( .A(rst), .B(Feedback[15]), .Z(
        PlaintextMUX_MUXInst_15_n2 ) );
  ORN2 PlaintextMUX_MUXInst_15_U1  ( .A(PlaintextMUX_MUXInst_15_n1 ), .B(
        PlaintextMUX_MUXInst_15_n2 ), .Z(StateRegInput[15]) );
  AND2 PlaintextMUX_MUXInst_16_U3  ( .A(Plaintext[16]), .B(rst), .Z(
        PlaintextMUX_MUXInst_16_n1 ) );
  ORN2 PlaintextMUX_MUXInst_16_U2  ( .A(rst), .B(Feedback[16]), .Z(
        PlaintextMUX_MUXInst_16_n2 ) );
  ORN2 PlaintextMUX_MUXInst_16_U1  ( .A(PlaintextMUX_MUXInst_16_n1 ), .B(
        PlaintextMUX_MUXInst_16_n2 ), .Z(StateRegInput[16]) );
  AND2 PlaintextMUX_MUXInst_17_U3  ( .A(Plaintext[17]), .B(rst), .Z(
        PlaintextMUX_MUXInst_17_n1 ) );
  ORN2 PlaintextMUX_MUXInst_17_U2  ( .A(rst), .B(Feedback[17]), .Z(
        PlaintextMUX_MUXInst_17_n2 ) );
  ORN2 PlaintextMUX_MUXInst_17_U1  ( .A(PlaintextMUX_MUXInst_17_n1 ), .B(
        PlaintextMUX_MUXInst_17_n2 ), .Z(StateRegInput[17]) );
  AND2 PlaintextMUX_MUXInst_18_U3  ( .A(Plaintext[18]), .B(rst), .Z(
        PlaintextMUX_MUXInst_18_n1 ) );
  ORN2 PlaintextMUX_MUXInst_18_U2  ( .A(rst), .B(Feedback[18]), .Z(
        PlaintextMUX_MUXInst_18_n2 ) );
  ORN2 PlaintextMUX_MUXInst_18_U1  ( .A(PlaintextMUX_MUXInst_18_n1 ), .B(
        PlaintextMUX_MUXInst_18_n2 ), .Z(StateRegInput[18]) );
  AND2 PlaintextMUX_MUXInst_19_U3  ( .A(Plaintext[19]), .B(rst), .Z(
        PlaintextMUX_MUXInst_19_n1 ) );
  ORN2 PlaintextMUX_MUXInst_19_U2  ( .A(rst), .B(Feedback[19]), .Z(
        PlaintextMUX_MUXInst_19_n2 ) );
  ORN2 PlaintextMUX_MUXInst_19_U1  ( .A(PlaintextMUX_MUXInst_19_n1 ), .B(
        PlaintextMUX_MUXInst_19_n2 ), .Z(StateRegInput[19]) );
  AND2 PlaintextMUX_MUXInst_20_U3  ( .A(Plaintext[20]), .B(rst), .Z(
        PlaintextMUX_MUXInst_20_n1 ) );
  ORN2 PlaintextMUX_MUXInst_20_U2  ( .A(rst), .B(Feedback[20]), .Z(
        PlaintextMUX_MUXInst_20_n2 ) );
  ORN2 PlaintextMUX_MUXInst_20_U1  ( .A(PlaintextMUX_MUXInst_20_n1 ), .B(
        PlaintextMUX_MUXInst_20_n2 ), .Z(StateRegInput[20]) );
  AND2 PlaintextMUX_MUXInst_21_U3  ( .A(Plaintext[21]), .B(rst), .Z(
        PlaintextMUX_MUXInst_21_n1 ) );
  ORN2 PlaintextMUX_MUXInst_21_U2  ( .A(rst), .B(Feedback[21]), .Z(
        PlaintextMUX_MUXInst_21_n2 ) );
  ORN2 PlaintextMUX_MUXInst_21_U1  ( .A(PlaintextMUX_MUXInst_21_n1 ), .B(
        PlaintextMUX_MUXInst_21_n2 ), .Z(StateRegInput[21]) );
  AND2 PlaintextMUX_MUXInst_22_U3  ( .A(Plaintext[22]), .B(rst), .Z(
        PlaintextMUX_MUXInst_22_n1 ) );
  ORN2 PlaintextMUX_MUXInst_22_U2  ( .A(rst), .B(Feedback[22]), .Z(
        PlaintextMUX_MUXInst_22_n2 ) );
  ORN2 PlaintextMUX_MUXInst_22_U1  ( .A(PlaintextMUX_MUXInst_22_n1 ), .B(
        PlaintextMUX_MUXInst_22_n2 ), .Z(StateRegInput[22]) );
  AND2 PlaintextMUX_MUXInst_23_U3  ( .A(Plaintext[23]), .B(rst), .Z(
        PlaintextMUX_MUXInst_23_n1 ) );
  ORN2 PlaintextMUX_MUXInst_23_U2  ( .A(rst), .B(Feedback[23]), .Z(
        PlaintextMUX_MUXInst_23_n2 ) );
  ORN2 PlaintextMUX_MUXInst_23_U1  ( .A(PlaintextMUX_MUXInst_23_n1 ), .B(
        PlaintextMUX_MUXInst_23_n2 ), .Z(StateRegInput[23]) );
  AND2 PlaintextMUX_MUXInst_24_U3  ( .A(Plaintext[24]), .B(rst), .Z(
        PlaintextMUX_MUXInst_24_n1 ) );
  ORN2 PlaintextMUX_MUXInst_24_U2  ( .A(rst), .B(Feedback[24]), .Z(
        PlaintextMUX_MUXInst_24_n2 ) );
  ORN2 PlaintextMUX_MUXInst_24_U1  ( .A(PlaintextMUX_MUXInst_24_n1 ), .B(
        PlaintextMUX_MUXInst_24_n2 ), .Z(StateRegInput[24]) );
  AND2 PlaintextMUX_MUXInst_25_U3  ( .A(Plaintext[25]), .B(rst), .Z(
        PlaintextMUX_MUXInst_25_n1 ) );
  ORN2 PlaintextMUX_MUXInst_25_U2  ( .A(rst), .B(Feedback[25]), .Z(
        PlaintextMUX_MUXInst_25_n2 ) );
  ORN2 PlaintextMUX_MUXInst_25_U1  ( .A(PlaintextMUX_MUXInst_25_n1 ), .B(
        PlaintextMUX_MUXInst_25_n2 ), .Z(StateRegInput[25]) );
  AND2 PlaintextMUX_MUXInst_26_U3  ( .A(Plaintext[26]), .B(rst), .Z(
        PlaintextMUX_MUXInst_26_n1 ) );
  ORN2 PlaintextMUX_MUXInst_26_U2  ( .A(rst), .B(Feedback[26]), .Z(
        PlaintextMUX_MUXInst_26_n2 ) );
  ORN2 PlaintextMUX_MUXInst_26_U1  ( .A(PlaintextMUX_MUXInst_26_n1 ), .B(
        PlaintextMUX_MUXInst_26_n2 ), .Z(StateRegInput[26]) );
  AND2 PlaintextMUX_MUXInst_27_U3  ( .A(Plaintext[27]), .B(rst), .Z(
        PlaintextMUX_MUXInst_27_n1 ) );
  ORN2 PlaintextMUX_MUXInst_27_U2  ( .A(rst), .B(Feedback[27]), .Z(
        PlaintextMUX_MUXInst_27_n2 ) );
  ORN2 PlaintextMUX_MUXInst_27_U1  ( .A(PlaintextMUX_MUXInst_27_n1 ), .B(
        PlaintextMUX_MUXInst_27_n2 ), .Z(StateRegInput[27]) );
  AND2 PlaintextMUX_MUXInst_28_U3  ( .A(Plaintext[28]), .B(rst), .Z(
        PlaintextMUX_MUXInst_28_n1 ) );
  ORN2 PlaintextMUX_MUXInst_28_U2  ( .A(rst), .B(Feedback[28]), .Z(
        PlaintextMUX_MUXInst_28_n2 ) );
  ORN2 PlaintextMUX_MUXInst_28_U1  ( .A(PlaintextMUX_MUXInst_28_n1 ), .B(
        PlaintextMUX_MUXInst_28_n2 ), .Z(StateRegInput[28]) );
  AND2 PlaintextMUX_MUXInst_29_U3  ( .A(Plaintext[29]), .B(rst), .Z(
        PlaintextMUX_MUXInst_29_n1 ) );
  ORN2 PlaintextMUX_MUXInst_29_U2  ( .A(rst), .B(Feedback[29]), .Z(
        PlaintextMUX_MUXInst_29_n2 ) );
  ORN2 PlaintextMUX_MUXInst_29_U1  ( .A(PlaintextMUX_MUXInst_29_n1 ), .B(
        PlaintextMUX_MUXInst_29_n2 ), .Z(StateRegInput[29]) );
  AND2 PlaintextMUX_MUXInst_30_U3  ( .A(Plaintext[30]), .B(rst), .Z(
        PlaintextMUX_MUXInst_30_n1 ) );
  ORN2 PlaintextMUX_MUXInst_30_U2  ( .A(rst), .B(Feedback[30]), .Z(
        PlaintextMUX_MUXInst_30_n2 ) );
  ORN2 PlaintextMUX_MUXInst_30_U1  ( .A(PlaintextMUX_MUXInst_30_n1 ), .B(
        PlaintextMUX_MUXInst_30_n2 ), .Z(StateRegInput[30]) );
  AND2 PlaintextMUX_MUXInst_31_U3  ( .A(Plaintext[31]), .B(rst), .Z(
        PlaintextMUX_MUXInst_31_n1 ) );
  ORN2 PlaintextMUX_MUXInst_31_U2  ( .A(rst), .B(Feedback[31]), .Z(
        PlaintextMUX_MUXInst_31_n2 ) );
  ORN2 PlaintextMUX_MUXInst_31_U1  ( .A(PlaintextMUX_MUXInst_31_n1 ), .B(
        PlaintextMUX_MUXInst_31_n2 ), .Z(StateRegInput[31]) );
  AND2 PlaintextMUX_MUXInst_32_U3  ( .A(Plaintext[32]), .B(rst), .Z(
        PlaintextMUX_MUXInst_32_n1 ) );
  ORN2 PlaintextMUX_MUXInst_32_U2  ( .A(rst), .B(Feedback[32]), .Z(
        PlaintextMUX_MUXInst_32_n2 ) );
  ORN2 PlaintextMUX_MUXInst_32_U1  ( .A(PlaintextMUX_MUXInst_32_n1 ), .B(
        PlaintextMUX_MUXInst_32_n2 ), .Z(StateRegInput[32]) );
  AND2 PlaintextMUX_MUXInst_33_U3  ( .A(Plaintext[33]), .B(rst), .Z(
        PlaintextMUX_MUXInst_33_n1 ) );
  ORN2 PlaintextMUX_MUXInst_33_U2  ( .A(rst), .B(Feedback[33]), .Z(
        PlaintextMUX_MUXInst_33_n2 ) );
  ORN2 PlaintextMUX_MUXInst_33_U1  ( .A(PlaintextMUX_MUXInst_33_n1 ), .B(
        PlaintextMUX_MUXInst_33_n2 ), .Z(StateRegInput[33]) );
  AND2 PlaintextMUX_MUXInst_34_U3  ( .A(Plaintext[34]), .B(rst), .Z(
        PlaintextMUX_MUXInst_34_n1 ) );
  ORN2 PlaintextMUX_MUXInst_34_U2  ( .A(rst), .B(Feedback[34]), .Z(
        PlaintextMUX_MUXInst_34_n2 ) );
  ORN2 PlaintextMUX_MUXInst_34_U1  ( .A(PlaintextMUX_MUXInst_34_n1 ), .B(
        PlaintextMUX_MUXInst_34_n2 ), .Z(StateRegInput[34]) );
  AND2 PlaintextMUX_MUXInst_35_U3  ( .A(Plaintext[35]), .B(rst), .Z(
        PlaintextMUX_MUXInst_35_n1 ) );
  ORN2 PlaintextMUX_MUXInst_35_U2  ( .A(rst), .B(Feedback[35]), .Z(
        PlaintextMUX_MUXInst_35_n2 ) );
  ORN2 PlaintextMUX_MUXInst_35_U1  ( .A(PlaintextMUX_MUXInst_35_n1 ), .B(
        PlaintextMUX_MUXInst_35_n2 ), .Z(StateRegInput[35]) );
  AND2 PlaintextMUX_MUXInst_36_U3  ( .A(Plaintext[36]), .B(rst), .Z(
        PlaintextMUX_MUXInst_36_n1 ) );
  ORN2 PlaintextMUX_MUXInst_36_U2  ( .A(rst), .B(Feedback[36]), .Z(
        PlaintextMUX_MUXInst_36_n2 ) );
  ORN2 PlaintextMUX_MUXInst_36_U1  ( .A(PlaintextMUX_MUXInst_36_n1 ), .B(
        PlaintextMUX_MUXInst_36_n2 ), .Z(StateRegInput[36]) );
  AND2 PlaintextMUX_MUXInst_37_U3  ( .A(Plaintext[37]), .B(rst), .Z(
        PlaintextMUX_MUXInst_37_n1 ) );
  ORN2 PlaintextMUX_MUXInst_37_U2  ( .A(rst), .B(Feedback[37]), .Z(
        PlaintextMUX_MUXInst_37_n2 ) );
  ORN2 PlaintextMUX_MUXInst_37_U1  ( .A(PlaintextMUX_MUXInst_37_n1 ), .B(
        PlaintextMUX_MUXInst_37_n2 ), .Z(StateRegInput[37]) );
  AND2 PlaintextMUX_MUXInst_38_U3  ( .A(Plaintext[38]), .B(rst), .Z(
        PlaintextMUX_MUXInst_38_n1 ) );
  ORN2 PlaintextMUX_MUXInst_38_U2  ( .A(rst), .B(Feedback[38]), .Z(
        PlaintextMUX_MUXInst_38_n2 ) );
  ORN2 PlaintextMUX_MUXInst_38_U1  ( .A(PlaintextMUX_MUXInst_38_n1 ), .B(
        PlaintextMUX_MUXInst_38_n2 ), .Z(StateRegInput[38]) );
  AND2 PlaintextMUX_MUXInst_39_U3  ( .A(Plaintext[39]), .B(rst), .Z(
        PlaintextMUX_MUXInst_39_n1 ) );
  ORN2 PlaintextMUX_MUXInst_39_U2  ( .A(rst), .B(Feedback[39]), .Z(
        PlaintextMUX_MUXInst_39_n2 ) );
  ORN2 PlaintextMUX_MUXInst_39_U1  ( .A(PlaintextMUX_MUXInst_39_n1 ), .B(
        PlaintextMUX_MUXInst_39_n2 ), .Z(StateRegInput[39]) );
  AND2 PlaintextMUX_MUXInst_40_U3  ( .A(Plaintext[40]), .B(rst), .Z(
        PlaintextMUX_MUXInst_40_n1 ) );
  ORN2 PlaintextMUX_MUXInst_40_U2  ( .A(rst), .B(Feedback[40]), .Z(
        PlaintextMUX_MUXInst_40_n2 ) );
  ORN2 PlaintextMUX_MUXInst_40_U1  ( .A(PlaintextMUX_MUXInst_40_n1 ), .B(
        PlaintextMUX_MUXInst_40_n2 ), .Z(StateRegInput[40]) );
  AND2 PlaintextMUX_MUXInst_41_U3  ( .A(Plaintext[41]), .B(rst), .Z(
        PlaintextMUX_MUXInst_41_n1 ) );
  ORN2 PlaintextMUX_MUXInst_41_U2  ( .A(rst), .B(Feedback[41]), .Z(
        PlaintextMUX_MUXInst_41_n2 ) );
  ORN2 PlaintextMUX_MUXInst_41_U1  ( .A(PlaintextMUX_MUXInst_41_n1 ), .B(
        PlaintextMUX_MUXInst_41_n2 ), .Z(StateRegInput[41]) );
  AND2 PlaintextMUX_MUXInst_42_U3  ( .A(Plaintext[42]), .B(rst), .Z(
        PlaintextMUX_MUXInst_42_n1 ) );
  ORN2 PlaintextMUX_MUXInst_42_U2  ( .A(rst), .B(Feedback[42]), .Z(
        PlaintextMUX_MUXInst_42_n2 ) );
  ORN2 PlaintextMUX_MUXInst_42_U1  ( .A(PlaintextMUX_MUXInst_42_n1 ), .B(
        PlaintextMUX_MUXInst_42_n2 ), .Z(StateRegInput[42]) );
  AND2 PlaintextMUX_MUXInst_43_U3  ( .A(Plaintext[43]), .B(rst), .Z(
        PlaintextMUX_MUXInst_43_n1 ) );
  ORN2 PlaintextMUX_MUXInst_43_U2  ( .A(rst), .B(Feedback[43]), .Z(
        PlaintextMUX_MUXInst_43_n2 ) );
  ORN2 PlaintextMUX_MUXInst_43_U1  ( .A(PlaintextMUX_MUXInst_43_n1 ), .B(
        PlaintextMUX_MUXInst_43_n2 ), .Z(StateRegInput[43]) );
  AND2 PlaintextMUX_MUXInst_44_U3  ( .A(Plaintext[44]), .B(rst), .Z(
        PlaintextMUX_MUXInst_44_n1 ) );
  ORN2 PlaintextMUX_MUXInst_44_U2  ( .A(rst), .B(Feedback[44]), .Z(
        PlaintextMUX_MUXInst_44_n2 ) );
  ORN2 PlaintextMUX_MUXInst_44_U1  ( .A(PlaintextMUX_MUXInst_44_n1 ), .B(
        PlaintextMUX_MUXInst_44_n2 ), .Z(StateRegInput[44]) );
  AND2 PlaintextMUX_MUXInst_45_U3  ( .A(Plaintext[45]), .B(rst), .Z(
        PlaintextMUX_MUXInst_45_n1 ) );
  ORN2 PlaintextMUX_MUXInst_45_U2  ( .A(rst), .B(Feedback[45]), .Z(
        PlaintextMUX_MUXInst_45_n2 ) );
  ORN2 PlaintextMUX_MUXInst_45_U1  ( .A(PlaintextMUX_MUXInst_45_n1 ), .B(
        PlaintextMUX_MUXInst_45_n2 ), .Z(StateRegInput[45]) );
  AND2 PlaintextMUX_MUXInst_46_U3  ( .A(Plaintext[46]), .B(rst), .Z(
        PlaintextMUX_MUXInst_46_n1 ) );
  ORN2 PlaintextMUX_MUXInst_46_U2  ( .A(rst), .B(Feedback[46]), .Z(
        PlaintextMUX_MUXInst_46_n2 ) );
  ORN2 PlaintextMUX_MUXInst_46_U1  ( .A(PlaintextMUX_MUXInst_46_n1 ), .B(
        PlaintextMUX_MUXInst_46_n2 ), .Z(StateRegInput[46]) );
  AND2 PlaintextMUX_MUXInst_47_U3  ( .A(Plaintext[47]), .B(rst), .Z(
        PlaintextMUX_MUXInst_47_n1 ) );
  ORN2 PlaintextMUX_MUXInst_47_U2  ( .A(rst), .B(Feedback[47]), .Z(
        PlaintextMUX_MUXInst_47_n2 ) );
  ORN2 PlaintextMUX_MUXInst_47_U1  ( .A(PlaintextMUX_MUXInst_47_n1 ), .B(
        PlaintextMUX_MUXInst_47_n2 ), .Z(StateRegInput[47]) );
  AND2 PlaintextMUX_MUXInst_48_U3  ( .A(Plaintext[48]), .B(rst), .Z(
        PlaintextMUX_MUXInst_48_n1 ) );
  ORN2 PlaintextMUX_MUXInst_48_U2  ( .A(rst), .B(Feedback[48]), .Z(
        PlaintextMUX_MUXInst_48_n2 ) );
  ORN2 PlaintextMUX_MUXInst_48_U1  ( .A(PlaintextMUX_MUXInst_48_n1 ), .B(
        PlaintextMUX_MUXInst_48_n2 ), .Z(StateRegInput[48]) );
  AND2 PlaintextMUX_MUXInst_49_U3  ( .A(Plaintext[49]), .B(rst), .Z(
        PlaintextMUX_MUXInst_49_n1 ) );
  ORN2 PlaintextMUX_MUXInst_49_U2  ( .A(rst), .B(Feedback[49]), .Z(
        PlaintextMUX_MUXInst_49_n2 ) );
  ORN2 PlaintextMUX_MUXInst_49_U1  ( .A(PlaintextMUX_MUXInst_49_n1 ), .B(
        PlaintextMUX_MUXInst_49_n2 ), .Z(StateRegInput[49]) );
  AND2 PlaintextMUX_MUXInst_50_U3  ( .A(Plaintext[50]), .B(rst), .Z(
        PlaintextMUX_MUXInst_50_n1 ) );
  ORN2 PlaintextMUX_MUXInst_50_U2  ( .A(rst), .B(Feedback[50]), .Z(
        PlaintextMUX_MUXInst_50_n2 ) );
  ORN2 PlaintextMUX_MUXInst_50_U1  ( .A(PlaintextMUX_MUXInst_50_n1 ), .B(
        PlaintextMUX_MUXInst_50_n2 ), .Z(StateRegInput[50]) );
  AND2 PlaintextMUX_MUXInst_51_U3  ( .A(Plaintext[51]), .B(rst), .Z(
        PlaintextMUX_MUXInst_51_n1 ) );
  ORN2 PlaintextMUX_MUXInst_51_U2  ( .A(rst), .B(Feedback[51]), .Z(
        PlaintextMUX_MUXInst_51_n2 ) );
  ORN2 PlaintextMUX_MUXInst_51_U1  ( .A(PlaintextMUX_MUXInst_51_n1 ), .B(
        PlaintextMUX_MUXInst_51_n2 ), .Z(StateRegInput[51]) );
  AND2 PlaintextMUX_MUXInst_52_U3  ( .A(Plaintext[52]), .B(rst), .Z(
        PlaintextMUX_MUXInst_52_n1 ) );
  ORN2 PlaintextMUX_MUXInst_52_U2  ( .A(rst), .B(Feedback[52]), .Z(
        PlaintextMUX_MUXInst_52_n2 ) );
  ORN2 PlaintextMUX_MUXInst_52_U1  ( .A(PlaintextMUX_MUXInst_52_n1 ), .B(
        PlaintextMUX_MUXInst_52_n2 ), .Z(StateRegInput[52]) );
  AND2 PlaintextMUX_MUXInst_53_U3  ( .A(Plaintext[53]), .B(rst), .Z(
        PlaintextMUX_MUXInst_53_n1 ) );
  ORN2 PlaintextMUX_MUXInst_53_U2  ( .A(rst), .B(Feedback[53]), .Z(
        PlaintextMUX_MUXInst_53_n2 ) );
  ORN2 PlaintextMUX_MUXInst_53_U1  ( .A(PlaintextMUX_MUXInst_53_n1 ), .B(
        PlaintextMUX_MUXInst_53_n2 ), .Z(StateRegInput[53]) );
  AND2 PlaintextMUX_MUXInst_54_U3  ( .A(Plaintext[54]), .B(rst), .Z(
        PlaintextMUX_MUXInst_54_n1 ) );
  ORN2 PlaintextMUX_MUXInst_54_U2  ( .A(rst), .B(Feedback[54]), .Z(
        PlaintextMUX_MUXInst_54_n2 ) );
  ORN2 PlaintextMUX_MUXInst_54_U1  ( .A(PlaintextMUX_MUXInst_54_n1 ), .B(
        PlaintextMUX_MUXInst_54_n2 ), .Z(StateRegInput[54]) );
  AND2 PlaintextMUX_MUXInst_55_U3  ( .A(Plaintext[55]), .B(rst), .Z(
        PlaintextMUX_MUXInst_55_n1 ) );
  ORN2 PlaintextMUX_MUXInst_55_U2  ( .A(rst), .B(Feedback[55]), .Z(
        PlaintextMUX_MUXInst_55_n2 ) );
  ORN2 PlaintextMUX_MUXInst_55_U1  ( .A(PlaintextMUX_MUXInst_55_n1 ), .B(
        PlaintextMUX_MUXInst_55_n2 ), .Z(StateRegInput[55]) );
  AND2 PlaintextMUX_MUXInst_56_U3  ( .A(Plaintext[56]), .B(rst), .Z(
        PlaintextMUX_MUXInst_56_n1 ) );
  ORN2 PlaintextMUX_MUXInst_56_U2  ( .A(rst), .B(Feedback[56]), .Z(
        PlaintextMUX_MUXInst_56_n2 ) );
  ORN2 PlaintextMUX_MUXInst_56_U1  ( .A(PlaintextMUX_MUXInst_56_n1 ), .B(
        PlaintextMUX_MUXInst_56_n2 ), .Z(StateRegInput[56]) );
  AND2 PlaintextMUX_MUXInst_57_U3  ( .A(Plaintext[57]), .B(rst), .Z(
        PlaintextMUX_MUXInst_57_n1 ) );
  ORN2 PlaintextMUX_MUXInst_57_U2  ( .A(rst), .B(Feedback[57]), .Z(
        PlaintextMUX_MUXInst_57_n2 ) );
  ORN2 PlaintextMUX_MUXInst_57_U1  ( .A(PlaintextMUX_MUXInst_57_n1 ), .B(
        PlaintextMUX_MUXInst_57_n2 ), .Z(StateRegInput[57]) );
  AND2 PlaintextMUX_MUXInst_58_U3  ( .A(Plaintext[58]), .B(rst), .Z(
        PlaintextMUX_MUXInst_58_n1 ) );
  ORN2 PlaintextMUX_MUXInst_58_U2  ( .A(rst), .B(Feedback[58]), .Z(
        PlaintextMUX_MUXInst_58_n2 ) );
  ORN2 PlaintextMUX_MUXInst_58_U1  ( .A(PlaintextMUX_MUXInst_58_n1 ), .B(
        PlaintextMUX_MUXInst_58_n2 ), .Z(StateRegInput[58]) );
  AND2 PlaintextMUX_MUXInst_59_U3  ( .A(Plaintext[59]), .B(rst), .Z(
        PlaintextMUX_MUXInst_59_n1 ) );
  ORN2 PlaintextMUX_MUXInst_59_U2  ( .A(rst), .B(Feedback[59]), .Z(
        PlaintextMUX_MUXInst_59_n2 ) );
  ORN2 PlaintextMUX_MUXInst_59_U1  ( .A(PlaintextMUX_MUXInst_59_n1 ), .B(
        PlaintextMUX_MUXInst_59_n2 ), .Z(StateRegInput[59]) );
  AND2 PlaintextMUX_MUXInst_60_U3  ( .A(Plaintext[60]), .B(rst), .Z(
        PlaintextMUX_MUXInst_60_n1 ) );
  ORN2 PlaintextMUX_MUXInst_60_U2  ( .A(rst), .B(Feedback[60]), .Z(
        PlaintextMUX_MUXInst_60_n2 ) );
  ORN2 PlaintextMUX_MUXInst_60_U1  ( .A(PlaintextMUX_MUXInst_60_n1 ), .B(
        PlaintextMUX_MUXInst_60_n2 ), .Z(StateRegInput[60]) );
  AND2 PlaintextMUX_MUXInst_61_U3  ( .A(Plaintext[61]), .B(rst), .Z(
        PlaintextMUX_MUXInst_61_n1 ) );
  ORN2 PlaintextMUX_MUXInst_61_U2  ( .A(rst), .B(Feedback[61]), .Z(
        PlaintextMUX_MUXInst_61_n2 ) );
  ORN2 PlaintextMUX_MUXInst_61_U1  ( .A(PlaintextMUX_MUXInst_61_n1 ), .B(
        PlaintextMUX_MUXInst_61_n2 ), .Z(StateRegInput[61]) );
  AND2 PlaintextMUX_MUXInst_62_U3  ( .A(Plaintext[62]), .B(rst), .Z(
        PlaintextMUX_MUXInst_62_n1 ) );
  ORN2 PlaintextMUX_MUXInst_62_U2  ( .A(rst), .B(Feedback[62]), .Z(
        PlaintextMUX_MUXInst_62_n2 ) );
  ORN2 PlaintextMUX_MUXInst_62_U1  ( .A(PlaintextMUX_MUXInst_62_n1 ), .B(
        PlaintextMUX_MUXInst_62_n2 ), .Z(StateRegInput[62]) );
  AND2 PlaintextMUX_MUXInst_63_U3  ( .A(Plaintext[63]), .B(rst), .Z(
        PlaintextMUX_MUXInst_63_n1 ) );
  ORN2 PlaintextMUX_MUXInst_63_U2  ( .A(rst), .B(Feedback[63]), .Z(
        PlaintextMUX_MUXInst_63_n2 ) );
  ORN2 PlaintextMUX_MUXInst_63_U1  ( .A(PlaintextMUX_MUXInst_63_n1 ), .B(
        PlaintextMUX_MUXInst_63_n2 ), .Z(StateRegInput[63]) );
  DFF StateReg_s_current_state_reg[0]  ( .D(StateRegInput[0]), .CP(clk), .Q(
        StateRegOutput[0]) );
  DFF StateReg_s_current_state_reg[1]  ( .D(StateRegInput[1]), .CP(clk), .Q(
        StateRegOutput[1]) );
  DFF StateReg_s_current_state_reg[2]  ( .D(StateRegInput[2]), .CP(clk), .Q(
        StateRegOutput[2]) );
  DFF StateReg_s_current_state_reg[3]  ( .D(StateRegInput[3]), .CP(clk), .Q(
        StateRegOutput[3]) );
  DFF StateReg_s_current_state_reg[4]  ( .D(StateRegInput[4]), .CP(clk), .Q(
        StateRegOutput[4]) );
  DFF StateReg_s_current_state_reg[5]  ( .D(StateRegInput[5]), .CP(clk), .Q(
        StateRegOutput[5]) );
  DFF StateReg_s_current_state_reg[6]  ( .D(StateRegInput[6]), .CP(clk), .Q(
        StateRegOutput[6]) );
  DFF StateReg_s_current_state_reg[7]  ( .D(StateRegInput[7]), .CP(clk), .Q(
        StateRegOutput[7]) );
  DFF StateReg_s_current_state_reg[8]  ( .D(StateRegInput[8]), .CP(clk), .Q(
        StateRegOutput[8]) );
  DFF StateReg_s_current_state_reg[9]  ( .D(StateRegInput[9]), .CP(clk), .Q(
        StateRegOutput[9]) );
  DFF StateReg_s_current_state_reg[10]  ( .D(StateRegInput[10]), .CP(clk), 
        .Q(StateRegOutput[10]) );
  DFF StateReg_s_current_state_reg[11]  ( .D(StateRegInput[11]), .CP(clk), 
        .Q(StateRegOutput[11]) );
  DFF StateReg_s_current_state_reg[12]  ( .D(StateRegInput[12]), .CP(clk), 
        .Q(StateRegOutput[12]) );
  DFF StateReg_s_current_state_reg[13]  ( .D(StateRegInput[13]), .CP(clk), 
        .Q(StateRegOutput[13]) );
  DFF StateReg_s_current_state_reg[14]  ( .D(StateRegInput[14]), .CP(clk), 
        .Q(StateRegOutput[14]) );
  DFF StateReg_s_current_state_reg[15]  ( .D(StateRegInput[15]), .CP(clk), 
        .Q(StateRegOutput[15]) );
  DFF StateReg_s_current_state_reg[16]  ( .D(StateRegInput[16]), .CP(clk), 
        .Q(StateRegOutput[16]) );
  DFF StateReg_s_current_state_reg[17]  ( .D(StateRegInput[17]), .CP(clk), 
        .Q(StateRegOutput[17]) );
  DFF StateReg_s_current_state_reg[18]  ( .D(StateRegInput[18]), .CP(clk), 
        .Q(StateRegOutput[18]) );
  DFF StateReg_s_current_state_reg[19]  ( .D(StateRegInput[19]), .CP(clk), 
        .Q(StateRegOutput[19]) );
  DFF StateReg_s_current_state_reg[20]  ( .D(StateRegInput[20]), .CP(clk), 
        .Q(StateRegOutput[20]) );
  DFF StateReg_s_current_state_reg[21]  ( .D(StateRegInput[21]), .CP(clk), 
        .Q(StateRegOutput[21]) );
  DFF StateReg_s_current_state_reg[22]  ( .D(StateRegInput[22]), .CP(clk), 
        .Q(StateRegOutput[22]) );
  DFF StateReg_s_current_state_reg[23]  ( .D(StateRegInput[23]), .CP(clk), 
        .Q(StateRegOutput[23]) );
  DFF StateReg_s_current_state_reg[24]  ( .D(StateRegInput[24]), .CP(clk), 
        .Q(StateRegOutput[24]) );
  DFF StateReg_s_current_state_reg[25]  ( .D(StateRegInput[25]), .CP(clk), 
        .Q(StateRegOutput[25]) );
  DFF StateReg_s_current_state_reg[26]  ( .D(StateRegInput[26]), .CP(clk), 
        .Q(StateRegOutput[26]) );
  DFF StateReg_s_current_state_reg[27]  ( .D(StateRegInput[27]), .CP(clk), 
        .Q(StateRegOutput[27]) );
  DFF StateReg_s_current_state_reg[28]  ( .D(StateRegInput[28]), .CP(clk), 
        .Q(StateRegOutput[28]) );
  DFF StateReg_s_current_state_reg[29]  ( .D(StateRegInput[29]), .CP(clk), 
        .Q(StateRegOutput[29]) );
  DFF StateReg_s_current_state_reg[30]  ( .D(StateRegInput[30]), .CP(clk), 
        .Q(StateRegOutput[30]) );
  DFF StateReg_s_current_state_reg[31]  ( .D(StateRegInput[31]), .CP(clk), 
        .Q(StateRegOutput[31]) );
  DFF StateReg_s_current_state_reg[32]  ( .D(StateRegInput[32]), .CP(clk), 
        .Q(StateRegOutput[32]) );
  DFF StateReg_s_current_state_reg[33]  ( .D(StateRegInput[33]), .CP(clk), 
        .Q(StateRegOutput[33]) );
  DFF StateReg_s_current_state_reg[34]  ( .D(StateRegInput[34]), .CP(clk), 
        .Q(StateRegOutput[34]) );
  DFF StateReg_s_current_state_reg[35]  ( .D(StateRegInput[35]), .CP(clk), 
        .Q(StateRegOutput[35]) );
  DFF StateReg_s_current_state_reg[36]  ( .D(StateRegInput[36]), .CP(clk), 
        .Q(StateRegOutput[36]) );
  DFF StateReg_s_current_state_reg[37]  ( .D(StateRegInput[37]), .CP(clk), 
        .Q(StateRegOutput[37]) );
  DFF StateReg_s_current_state_reg[38]  ( .D(StateRegInput[38]), .CP(clk), 
        .Q(StateRegOutput[38]) );
  DFF StateReg_s_current_state_reg[39]  ( .D(StateRegInput[39]), .CP(clk), 
        .Q(StateRegOutput[39]) );
  DFF StateReg_s_current_state_reg[40]  ( .D(StateRegInput[40]), .CP(clk), 
        .Q(StateRegOutput[40]) );
  DFF StateReg_s_current_state_reg[41]  ( .D(StateRegInput[41]), .CP(clk), 
        .Q(StateRegOutput[41]) );
  DFF StateReg_s_current_state_reg[42]  ( .D(StateRegInput[42]), .CP(clk), 
        .Q(StateRegOutput[42]) );
  DFF StateReg_s_current_state_reg[43]  ( .D(StateRegInput[43]), .CP(clk), 
        .Q(StateRegOutput[43]) );
  DFF StateReg_s_current_state_reg[44]  ( .D(StateRegInput[44]), .CP(clk), 
        .Q(StateRegOutput[44]) );
  DFF StateReg_s_current_state_reg[45]  ( .D(StateRegInput[45]), .CP(clk), 
        .Q(StateRegOutput[45]) );
  DFF StateReg_s_current_state_reg[46]  ( .D(StateRegInput[46]), .CP(clk), 
        .Q(StateRegOutput[46]) );
  DFF StateReg_s_current_state_reg[47]  ( .D(StateRegInput[47]), .CP(clk), 
        .Q(StateRegOutput[47]) );
  DFF StateReg_s_current_state_reg[48]  ( .D(StateRegInput[48]), .CP(clk), 
        .Q(StateRegOutput[48]) );
  DFF StateReg_s_current_state_reg[49]  ( .D(StateRegInput[49]), .CP(clk), 
        .Q(StateRegOutput[49]) );
  DFF StateReg_s_current_state_reg[50]  ( .D(StateRegInput[50]), .CP(clk), 
        .Q(StateRegOutput[50]) );
  DFF StateReg_s_current_state_reg[51]  ( .D(StateRegInput[51]), .CP(clk), 
        .Q(StateRegOutput[51]) );
  DFF StateReg_s_current_state_reg[52]  ( .D(StateRegInput[52]), .CP(clk), 
        .Q(StateRegOutput[52]) );
  DFF StateReg_s_current_state_reg[53]  ( .D(StateRegInput[53]), .CP(clk), 
        .Q(StateRegOutput[53]) );
  DFF StateReg_s_current_state_reg[54]  ( .D(StateRegInput[54]), .CP(clk), 
        .Q(StateRegOutput[54]) );
  DFF StateReg_s_current_state_reg[55]  ( .D(StateRegInput[55]), .CP(clk), 
        .Q(StateRegOutput[55]) );
  DFF StateReg_s_current_state_reg[56]  ( .D(StateRegInput[56]), .CP(clk), 
        .Q(StateRegOutput[56]) );
  DFF StateReg_s_current_state_reg[57]  ( .D(StateRegInput[57]), .CP(clk), 
        .Q(StateRegOutput[57]) );
  DFF StateReg_s_current_state_reg[58]  ( .D(StateRegInput[58]), .CP(clk), 
        .Q(StateRegOutput[58]) );
  DFF StateReg_s_current_state_reg[59]  ( .D(StateRegInput[59]), .CP(clk), 
        .Q(StateRegOutput[59]) );
  DFF StateReg_s_current_state_reg[60]  ( .D(StateRegInput[60]), .CP(clk), 
        .Q(StateRegOutput[60]) );
  DFF StateReg_s_current_state_reg[61]  ( .D(StateRegInput[61]), .CP(clk), 
        .Q(StateRegOutput[61]) );
  DFF StateReg_s_current_state_reg[62]  ( .D(StateRegInput[62]), .CP(clk), 
        .Q(StateRegOutput[62]) );
  DFF StateReg_s_current_state_reg[63]  ( .D(StateRegInput[63]), .CP(clk), 
        .Q(StateRegOutput[63]) );
  XOR2 AddKeyXOR_XORInst_0_0_U2  ( .A(Key[0]), .B(StateRegOutput[0]), .Z(
        AddKeyXOR_XORInst_0_0_n1 ) );
  XOR2 AddKeyXOR_XORInst_0_0_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_0_0_n1 ), 
        .Z(Ciphertext[0]) );
  XOR2 AddKeyXOR_XORInst_0_1_U2  ( .A(Key[1]), .B(StateRegOutput[1]), .Z(
        AddKeyXOR_XORInst_0_1_n1 ) );
  XOR2 AddKeyXOR_XORInst_0_1_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_0_1_n1 ), 
        .Z(Ciphertext[1]) );
  XOR2 AddKeyXOR_XORInst_0_2_U2  ( .A(Key[2]), .B(StateRegOutput[2]), .Z(
        AddKeyXOR_XORInst_0_2_n1 ) );
  XOR2 AddKeyXOR_XORInst_0_2_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_0_2_n1 ), 
        .Z(Ciphertext[2]) );
  XOR2 AddKeyXOR_XORInst_0_3_U2  ( .A(Key[3]), .B(StateRegOutput[3]), .Z(
        AddKeyXOR_XORInst_0_3_n1 ) );
  XOR2 AddKeyXOR_XORInst_0_3_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_0_3_n1 ), 
        .Z(Ciphertext[3]) );
  XOR2 AddKeyXOR_XORInst_1_0_U2  ( .A(Key[4]), .B(StateRegOutput[4]), .Z(
        AddKeyXOR_XORInst_1_0_n1 ) );
  XOR2 AddKeyXOR_XORInst_1_0_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_1_0_n1 ), 
        .Z(Ciphertext[4]) );
  XOR2 AddKeyXOR_XORInst_1_1_U2  ( .A(Key[5]), .B(StateRegOutput[5]), .Z(
        AddKeyXOR_XORInst_1_1_n1 ) );
  XOR2 AddKeyXOR_XORInst_1_1_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_1_1_n1 ), 
        .Z(Ciphertext[5]) );
  XOR2 AddKeyXOR_XORInst_1_2_U2  ( .A(Key[6]), .B(StateRegOutput[6]), .Z(
        AddKeyXOR_XORInst_1_2_n1 ) );
  XOR2 AddKeyXOR_XORInst_1_2_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_1_2_n1 ), 
        .Z(Ciphertext[6]) );
  XOR2 AddKeyXOR_XORInst_1_3_U2  ( .A(Key[7]), .B(StateRegOutput[7]), .Z(
        AddKeyXOR_XORInst_1_3_n1 ) );
  XOR2 AddKeyXOR_XORInst_1_3_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_1_3_n1 ), 
        .Z(Ciphertext[7]) );
  XOR2 AddKeyXOR_XORInst_2_0_U2  ( .A(Key[8]), .B(StateRegOutput[8]), .Z(
        AddKeyXOR_XORInst_2_0_n1 ) );
  XOR2 AddKeyXOR_XORInst_2_0_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_2_0_n1 ), 
        .Z(Ciphertext[8]) );
  XOR2 AddKeyXOR_XORInst_2_1_U2  ( .A(Key[9]), .B(StateRegOutput[9]), .Z(
        AddKeyXOR_XORInst_2_1_n1 ) );
  XOR2 AddKeyXOR_XORInst_2_1_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_2_1_n1 ), 
        .Z(Ciphertext[9]) );
  XOR2 AddKeyXOR_XORInst_2_2_U2  ( .A(Key[10]), .B(StateRegOutput[10]), .Z(
        AddKeyXOR_XORInst_2_2_n1 ) );
  XOR2 AddKeyXOR_XORInst_2_2_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_2_2_n1 ), 
        .Z(Ciphertext[10]) );
  XOR2 AddKeyXOR_XORInst_2_3_U2  ( .A(Key[11]), .B(StateRegOutput[11]), .Z(
        AddKeyXOR_XORInst_2_3_n1 ) );
  XOR2 AddKeyXOR_XORInst_2_3_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_2_3_n1 ), 
        .Z(Ciphertext[11]) );
  XOR2 AddKeyXOR_XORInst_3_0_U2  ( .A(Key[12]), .B(StateRegOutput[12]), .Z(
        AddKeyXOR_XORInst_3_0_n1 ) );
  XOR2 AddKeyXOR_XORInst_3_0_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_3_0_n1 ), 
        .Z(Ciphertext[12]) );
  XOR2 AddKeyXOR_XORInst_3_1_U2  ( .A(Key[13]), .B(StateRegOutput[13]), .Z(
        AddKeyXOR_XORInst_3_1_n1 ) );
  XOR2 AddKeyXOR_XORInst_3_1_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_3_1_n1 ), 
        .Z(Ciphertext[13]) );
  XOR2 AddKeyXOR_XORInst_3_2_U2  ( .A(Key[14]), .B(StateRegOutput[14]), .Z(
        AddKeyXOR_XORInst_3_2_n1 ) );
  XOR2 AddKeyXOR_XORInst_3_2_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_3_2_n1 ), 
        .Z(Ciphertext[14]) );
  XOR2 AddKeyXOR_XORInst_3_3_U2  ( .A(Key[15]), .B(StateRegOutput[15]), .Z(
        AddKeyXOR_XORInst_3_3_n1 ) );
  XOR2 AddKeyXOR_XORInst_3_3_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_3_3_n1 ), 
        .Z(Ciphertext[15]) );
  XOR2 AddKeyXOR_XORInst_4_0_U2  ( .A(Key[16]), .B(StateRegOutput[16]), .Z(
        AddKeyXOR_XORInst_4_0_n1 ) );
  XOR2 AddKeyXOR_XORInst_4_0_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_4_0_n1 ), 
        .Z(Ciphertext[16]) );
  XOR2 AddKeyXOR_XORInst_4_1_U2  ( .A(Key[17]), .B(StateRegOutput[17]), .Z(
        AddKeyXOR_XORInst_4_1_n1 ) );
  XOR2 AddKeyXOR_XORInst_4_1_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_4_1_n1 ), 
        .Z(Ciphertext[17]) );
  XOR2 AddKeyXOR_XORInst_4_2_U2  ( .A(Key[18]), .B(StateRegOutput[18]), .Z(
        AddKeyXOR_XORInst_4_2_n1 ) );
  XOR2 AddKeyXOR_XORInst_4_2_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_4_2_n1 ), 
        .Z(Ciphertext[18]) );
  XOR2 AddKeyXOR_XORInst_4_3_U2  ( .A(Key[19]), .B(StateRegOutput[19]), .Z(
        AddKeyXOR_XORInst_4_3_n1 ) );
  XOR2 AddKeyXOR_XORInst_4_3_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_4_3_n1 ), 
        .Z(Ciphertext[19]) );
  XOR2 AddKeyXOR_XORInst_5_0_U2  ( .A(Key[20]), .B(StateRegOutput[20]), .Z(
        AddKeyXOR_XORInst_5_0_n1 ) );
  XOR2 AddKeyXOR_XORInst_5_0_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_5_0_n1 ), 
        .Z(Ciphertext[20]) );
  XOR2 AddKeyXOR_XORInst_5_1_U2  ( .A(Key[21]), .B(StateRegOutput[21]), .Z(
        AddKeyXOR_XORInst_5_1_n1 ) );
  XOR2 AddKeyXOR_XORInst_5_1_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_5_1_n1 ), 
        .Z(Ciphertext[21]) );
  XOR2 AddKeyXOR_XORInst_5_2_U2  ( .A(Key[22]), .B(StateRegOutput[22]), .Z(
        AddKeyXOR_XORInst_5_2_n1 ) );
  XOR2 AddKeyXOR_XORInst_5_2_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_5_2_n1 ), 
        .Z(Ciphertext[22]) );
  XOR2 AddKeyXOR_XORInst_5_3_U2  ( .A(Key[23]), .B(StateRegOutput[23]), .Z(
        AddKeyXOR_XORInst_5_3_n1 ) );
  XOR2 AddKeyXOR_XORInst_5_3_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_5_3_n1 ), 
        .Z(Ciphertext[23]) );
  XOR2 AddKeyXOR_XORInst_6_0_U2  ( .A(Key[24]), .B(StateRegOutput[24]), .Z(
        AddKeyXOR_XORInst_6_0_n1 ) );
  XOR2 AddKeyXOR_XORInst_6_0_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_6_0_n1 ), 
        .Z(Ciphertext[24]) );
  XOR2 AddKeyXOR_XORInst_6_1_U2  ( .A(Key[25]), .B(StateRegOutput[25]), .Z(
        AddKeyXOR_XORInst_6_1_n1 ) );
  XOR2 AddKeyXOR_XORInst_6_1_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_6_1_n1 ), 
        .Z(Ciphertext[25]) );
  XOR2 AddKeyXOR_XORInst_6_2_U2  ( .A(Key[26]), .B(StateRegOutput[26]), .Z(
        AddKeyXOR_XORInst_6_2_n1 ) );
  XOR2 AddKeyXOR_XORInst_6_2_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_6_2_n1 ), 
        .Z(Ciphertext[26]) );
  XOR2 AddKeyXOR_XORInst_6_3_U2  ( .A(Key[27]), .B(StateRegOutput[27]), .Z(
        AddKeyXOR_XORInst_6_3_n1 ) );
  XOR2 AddKeyXOR_XORInst_6_3_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_6_3_n1 ), 
        .Z(Ciphertext[27]) );
  XOR2 AddKeyXOR_XORInst_7_0_U2  ( .A(Key[28]), .B(StateRegOutput[28]), .Z(
        AddKeyXOR_XORInst_7_0_n1 ) );
  XOR2 AddKeyXOR_XORInst_7_0_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_7_0_n1 ), 
        .Z(Ciphertext[28]) );
  XOR2 AddKeyXOR_XORInst_7_1_U2  ( .A(Key[29]), .B(StateRegOutput[29]), .Z(
        AddKeyXOR_XORInst_7_1_n1 ) );
  XOR2 AddKeyXOR_XORInst_7_1_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_7_1_n1 ), 
        .Z(Ciphertext[29]) );
  XOR2 AddKeyXOR_XORInst_7_2_U2  ( .A(Key[30]), .B(StateRegOutput[30]), .Z(
        AddKeyXOR_XORInst_7_2_n1 ) );
  XOR2 AddKeyXOR_XORInst_7_2_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_7_2_n1 ), 
        .Z(Ciphertext[30]) );
  XOR2 AddKeyXOR_XORInst_7_3_U2  ( .A(Key[31]), .B(StateRegOutput[31]), .Z(
        AddKeyXOR_XORInst_7_3_n1 ) );
  XOR2 AddKeyXOR_XORInst_7_3_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_7_3_n1 ), 
        .Z(Ciphertext[31]) );
  XOR2 AddKeyXOR_XORInst_8_0_U2  ( .A(Key[32]), .B(StateRegOutput[32]), .Z(
        AddKeyXOR_XORInst_8_0_n1 ) );
  XOR2 AddKeyXOR_XORInst_8_0_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_8_0_n1 ), 
        .Z(Ciphertext[32]) );
  XOR2 AddKeyXOR_XORInst_8_1_U2  ( .A(Key[33]), .B(StateRegOutput[33]), .Z(
        AddKeyXOR_XORInst_8_1_n1 ) );
  XOR2 AddKeyXOR_XORInst_8_1_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_8_1_n1 ), 
        .Z(Ciphertext[33]) );
  XOR2 AddKeyXOR_XORInst_8_2_U2  ( .A(Key[34]), .B(StateRegOutput[34]), .Z(
        AddKeyXOR_XORInst_8_2_n1 ) );
  XOR2 AddKeyXOR_XORInst_8_2_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_8_2_n1 ), 
        .Z(Ciphertext[34]) );
  XOR2 AddKeyXOR_XORInst_8_3_U2  ( .A(Key[35]), .B(StateRegOutput[35]), .Z(
        AddKeyXOR_XORInst_8_3_n1 ) );
  XOR2 AddKeyXOR_XORInst_8_3_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_8_3_n1 ), 
        .Z(Ciphertext[35]) );
  XOR2 AddKeyXOR_XORInst_9_0_U2  ( .A(Key[36]), .B(StateRegOutput[36]), .Z(
        AddKeyXOR_XORInst_9_0_n1 ) );
  XOR2 AddKeyXOR_XORInst_9_0_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_9_0_n1 ), 
        .Z(Ciphertext[36]) );
  XOR2 AddKeyXOR_XORInst_9_1_U2  ( .A(Key[37]), .B(StateRegOutput[37]), .Z(
        AddKeyXOR_XORInst_9_1_n1 ) );
  XOR2 AddKeyXOR_XORInst_9_1_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_9_1_n1 ), 
        .Z(Ciphertext[37]) );
  XOR2 AddKeyXOR_XORInst_9_2_U2  ( .A(Key[38]), .B(StateRegOutput[38]), .Z(
        AddKeyXOR_XORInst_9_2_n1 ) );
  XOR2 AddKeyXOR_XORInst_9_2_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_9_2_n1 ), 
        .Z(Ciphertext[38]) );
  XOR2 AddKeyXOR_XORInst_9_3_U2  ( .A(Key[39]), .B(StateRegOutput[39]), .Z(
        AddKeyXOR_XORInst_9_3_n1 ) );
  XOR2 AddKeyXOR_XORInst_9_3_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_9_3_n1 ), 
        .Z(Ciphertext[39]) );
  XOR2 AddKeyXOR_XORInst_10_0_U2  ( .A(Key[40]), .B(StateRegOutput[40]), .Z(
        AddKeyXOR_XORInst_10_0_n1 ) );
  XOR2 AddKeyXOR_XORInst_10_0_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_10_0_n1 ), 
        .Z(Ciphertext[40]) );
  XOR2 AddKeyXOR_XORInst_10_1_U2  ( .A(Key[41]), .B(StateRegOutput[41]), .Z(
        AddKeyXOR_XORInst_10_1_n1 ) );
  XOR2 AddKeyXOR_XORInst_10_1_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_10_1_n1 ), 
        .Z(Ciphertext[41]) );
  XOR2 AddKeyXOR_XORInst_10_2_U2  ( .A(Key[42]), .B(StateRegOutput[42]), .Z(
        AddKeyXOR_XORInst_10_2_n1 ) );
  XOR2 AddKeyXOR_XORInst_10_2_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_10_2_n1 ), 
        .Z(Ciphertext[42]) );
  XOR2 AddKeyXOR_XORInst_10_3_U2  ( .A(Key[43]), .B(StateRegOutput[43]), .Z(
        AddKeyXOR_XORInst_10_3_n1 ) );
  XOR2 AddKeyXOR_XORInst_10_3_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_10_3_n1 ), 
        .Z(Ciphertext[43]) );
  XOR2 AddKeyXOR_XORInst_11_0_U2  ( .A(Key[44]), .B(StateRegOutput[44]), .Z(
        AddKeyXOR_XORInst_11_0_n1 ) );
  XOR2 AddKeyXOR_XORInst_11_0_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_11_0_n1 ), 
        .Z(Ciphertext[44]) );
  XOR2 AddKeyXOR_XORInst_11_1_U2  ( .A(Key[45]), .B(StateRegOutput[45]), .Z(
        AddKeyXOR_XORInst_11_1_n1 ) );
  XOR2 AddKeyXOR_XORInst_11_1_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_11_1_n1 ), 
        .Z(Ciphertext[45]) );
  XOR2 AddKeyXOR_XORInst_11_2_U2  ( .A(Key[46]), .B(StateRegOutput[46]), .Z(
        AddKeyXOR_XORInst_11_2_n1 ) );
  XOR2 AddKeyXOR_XORInst_11_2_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_11_2_n1 ), 
        .Z(Ciphertext[46]) );
  XOR2 AddKeyXOR_XORInst_11_3_U2  ( .A(Key[47]), .B(StateRegOutput[47]), .Z(
        AddKeyXOR_XORInst_11_3_n1 ) );
  XOR2 AddKeyXOR_XORInst_11_3_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_11_3_n1 ), 
        .Z(Ciphertext[47]) );
  XOR2 AddKeyXOR_XORInst_12_0_U2  ( .A(Key[48]), .B(StateRegOutput[48]), .Z(
        AddKeyXOR_XORInst_12_0_n1 ) );
  XOR2 AddKeyXOR_XORInst_12_0_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_12_0_n1 ), 
        .Z(Ciphertext[48]) );
  XOR2 AddKeyXOR_XORInst_12_1_U2  ( .A(Key[49]), .B(StateRegOutput[49]), .Z(
        AddKeyXOR_XORInst_12_1_n1 ) );
  XOR2 AddKeyXOR_XORInst_12_1_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_12_1_n1 ), 
        .Z(Ciphertext[49]) );
  XOR2 AddKeyXOR_XORInst_12_2_U2  ( .A(Key[50]), .B(StateRegOutput[50]), .Z(
        AddKeyXOR_XORInst_12_2_n1 ) );
  XOR2 AddKeyXOR_XORInst_12_2_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_12_2_n1 ), 
        .Z(Ciphertext[50]) );
  XOR2 AddKeyXOR_XORInst_12_3_U2  ( .A(Key[51]), .B(StateRegOutput[51]), .Z(
        AddKeyXOR_XORInst_12_3_n1 ) );
  XOR2 AddKeyXOR_XORInst_12_3_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_12_3_n1 ), 
        .Z(Ciphertext[51]) );
  XOR2 AddKeyXOR_XORInst_13_0_U2  ( .A(Key[52]), .B(StateRegOutput[52]), .Z(
        AddKeyXOR_XORInst_13_0_n1 ) );
  XOR2 AddKeyXOR_XORInst_13_0_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_13_0_n1 ), 
        .Z(Ciphertext[52]) );
  XOR2 AddKeyXOR_XORInst_13_1_U2  ( .A(Key[53]), .B(StateRegOutput[53]), .Z(
        AddKeyXOR_XORInst_13_1_n1 ) );
  XOR2 AddKeyXOR_XORInst_13_1_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_13_1_n1 ), 
        .Z(Ciphertext[53]) );
  XOR2 AddKeyXOR_XORInst_13_2_U2  ( .A(Key[54]), .B(StateRegOutput[54]), .Z(
        AddKeyXOR_XORInst_13_2_n1 ) );
  XOR2 AddKeyXOR_XORInst_13_2_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_13_2_n1 ), 
        .Z(Ciphertext[54]) );
  XOR2 AddKeyXOR_XORInst_13_3_U2  ( .A(Key[55]), .B(StateRegOutput[55]), .Z(
        AddKeyXOR_XORInst_13_3_n1 ) );
  XOR2 AddKeyXOR_XORInst_13_3_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_13_3_n1 ), 
        .Z(Ciphertext[55]) );
  XOR2 AddKeyXOR_XORInst_14_0_U2  ( .A(Key[56]), .B(StateRegOutput[56]), .Z(
        AddKeyXOR_XORInst_14_0_n1 ) );
  XOR2 AddKeyXOR_XORInst_14_0_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_14_0_n1 ), 
        .Z(Ciphertext[56]) );
  XOR2 AddKeyXOR_XORInst_14_1_U2  ( .A(Key[57]), .B(StateRegOutput[57]), .Z(
        AddKeyXOR_XORInst_14_1_n1 ) );
  XOR2 AddKeyXOR_XORInst_14_1_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_14_1_n1 ), 
        .Z(Ciphertext[57]) );
  XOR2 AddKeyXOR_XORInst_14_2_U2  ( .A(Key[58]), .B(StateRegOutput[58]), .Z(
        AddKeyXOR_XORInst_14_2_n1 ) );
  XOR2 AddKeyXOR_XORInst_14_2_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_14_2_n1 ), 
        .Z(Ciphertext[58]) );
  XOR2 AddKeyXOR_XORInst_14_3_U2  ( .A(Key[59]), .B(StateRegOutput[59]), .Z(
        AddKeyXOR_XORInst_14_3_n1 ) );
  XOR2 AddKeyXOR_XORInst_14_3_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_14_3_n1 ), 
        .Z(Ciphertext[59]) );
  XOR2 AddKeyXOR_XORInst_15_0_U2  ( .A(Key[60]), .B(StateRegOutput[60]), .Z(
        AddKeyXOR_XORInst_15_0_n1 ) );
  XOR2 AddKeyXOR_XORInst_15_0_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_15_0_n1 ), 
        .Z(Ciphertext[60]) );
  XOR2 AddKeyXOR_XORInst_15_1_U2  ( .A(Key[61]), .B(StateRegOutput[61]), .Z(
        AddKeyXOR_XORInst_15_1_n1 ) );
  XOR2 AddKeyXOR_XORInst_15_1_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_15_1_n1 ), 
        .Z(Ciphertext[61]) );
  XOR2 AddKeyXOR_XORInst_15_2_U2  ( .A(Key[62]), .B(StateRegOutput[62]), .Z(
        AddKeyXOR_XORInst_15_2_n1 ) );
  XOR2 AddKeyXOR_XORInst_15_2_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_15_2_n1 ), 
        .Z(Ciphertext[62]) );
  XOR2 AddKeyXOR_XORInst_15_3_U2  ( .A(Key[63]), .B(StateRegOutput[63]), .Z(
        AddKeyXOR_XORInst_15_3_n1 ) );
  XOR2 AddKeyXOR_XORInst_15_3_U1  ( .A(1'b0), .B(AddKeyXOR_XORInst_15_3_n1 ), 
        .Z(Ciphertext[63]) );
  AND2 AddKeyMUX_MUXInst_0_U3  ( .A(Ciphertext[0]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_0_n1 ) );
  ORN2 AddKeyMUX_MUXInst_0_U2  ( .A(AddKey), .B(StateRegOutput[0]), .Z(
        AddKeyMUX_MUXInst_0_n2 ) );
  ORN2 AddKeyMUX_MUXInst_0_U1  ( .A(AddKeyMUX_MUXInst_0_n1 ), .B(
        AddKeyMUX_MUXInst_0_n2 ), .Z(AddKeyMUXOutput[0]) );
  AND2 AddKeyMUX_MUXInst_1_U3  ( .A(Ciphertext[1]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_1_n1 ) );
  ORN2 AddKeyMUX_MUXInst_1_U2  ( .A(AddKey), .B(StateRegOutput[1]), .Z(
        AddKeyMUX_MUXInst_1_n2 ) );
  ORN2 AddKeyMUX_MUXInst_1_U1  ( .A(AddKeyMUX_MUXInst_1_n1 ), .B(
        AddKeyMUX_MUXInst_1_n2 ), .Z(AddKeyMUXOutput[1]) );
  AND2 AddKeyMUX_MUXInst_2_U3  ( .A(Ciphertext[2]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_2_n1 ) );
  ORN2 AddKeyMUX_MUXInst_2_U2  ( .A(AddKey), .B(StateRegOutput[2]), .Z(
        AddKeyMUX_MUXInst_2_n2 ) );
  ORN2 AddKeyMUX_MUXInst_2_U1  ( .A(AddKeyMUX_MUXInst_2_n1 ), .B(
        AddKeyMUX_MUXInst_2_n2 ), .Z(AddKeyMUXOutput[2]) );
  AND2 AddKeyMUX_MUXInst_3_U3  ( .A(Ciphertext[3]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_3_n1 ) );
  ORN2 AddKeyMUX_MUXInst_3_U2  ( .A(AddKey), .B(StateRegOutput[3]), .Z(
        AddKeyMUX_MUXInst_3_n2 ) );
  ORN2 AddKeyMUX_MUXInst_3_U1  ( .A(AddKeyMUX_MUXInst_3_n1 ), .B(
        AddKeyMUX_MUXInst_3_n2 ), .Z(AddKeyMUXOutput[3]) );
  AND2 AddKeyMUX_MUXInst_4_U3  ( .A(Ciphertext[4]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_4_n1 ) );
  ORN2 AddKeyMUX_MUXInst_4_U2  ( .A(AddKey), .B(StateRegOutput[4]), .Z(
        AddKeyMUX_MUXInst_4_n2 ) );
  ORN2 AddKeyMUX_MUXInst_4_U1  ( .A(AddKeyMUX_MUXInst_4_n1 ), .B(
        AddKeyMUX_MUXInst_4_n2 ), .Z(AddKeyMUXOutput[4]) );
  AND2 AddKeyMUX_MUXInst_5_U3  ( .A(Ciphertext[5]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_5_n1 ) );
  ORN2 AddKeyMUX_MUXInst_5_U2  ( .A(AddKey), .B(StateRegOutput[5]), .Z(
        AddKeyMUX_MUXInst_5_n2 ) );
  ORN2 AddKeyMUX_MUXInst_5_U1  ( .A(AddKeyMUX_MUXInst_5_n1 ), .B(
        AddKeyMUX_MUXInst_5_n2 ), .Z(AddKeyMUXOutput[5]) );
  AND2 AddKeyMUX_MUXInst_6_U3  ( .A(Ciphertext[6]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_6_n1 ) );
  ORN2 AddKeyMUX_MUXInst_6_U2  ( .A(AddKey), .B(StateRegOutput[6]), .Z(
        AddKeyMUX_MUXInst_6_n2 ) );
  ORN2 AddKeyMUX_MUXInst_6_U1  ( .A(AddKeyMUX_MUXInst_6_n1 ), .B(
        AddKeyMUX_MUXInst_6_n2 ), .Z(AddKeyMUXOutput[6]) );
  AND2 AddKeyMUX_MUXInst_7_U3  ( .A(Ciphertext[7]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_7_n1 ) );
  ORN2 AddKeyMUX_MUXInst_7_U2  ( .A(AddKey), .B(StateRegOutput[7]), .Z(
        AddKeyMUX_MUXInst_7_n2 ) );
  ORN2 AddKeyMUX_MUXInst_7_U1  ( .A(AddKeyMUX_MUXInst_7_n1 ), .B(
        AddKeyMUX_MUXInst_7_n2 ), .Z(AddKeyMUXOutput[7]) );
  AND2 AddKeyMUX_MUXInst_8_U3  ( .A(Ciphertext[8]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_8_n1 ) );
  ORN2 AddKeyMUX_MUXInst_8_U2  ( .A(AddKey), .B(StateRegOutput[8]), .Z(
        AddKeyMUX_MUXInst_8_n2 ) );
  ORN2 AddKeyMUX_MUXInst_8_U1  ( .A(AddKeyMUX_MUXInst_8_n1 ), .B(
        AddKeyMUX_MUXInst_8_n2 ), .Z(AddKeyMUXOutput[8]) );
  AND2 AddKeyMUX_MUXInst_9_U3  ( .A(Ciphertext[9]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_9_n1 ) );
  ORN2 AddKeyMUX_MUXInst_9_U2  ( .A(AddKey), .B(StateRegOutput[9]), .Z(
        AddKeyMUX_MUXInst_9_n2 ) );
  ORN2 AddKeyMUX_MUXInst_9_U1  ( .A(AddKeyMUX_MUXInst_9_n1 ), .B(
        AddKeyMUX_MUXInst_9_n2 ), .Z(AddKeyMUXOutput[9]) );
  AND2 AddKeyMUX_MUXInst_10_U3  ( .A(Ciphertext[10]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_10_n1 ) );
  ORN2 AddKeyMUX_MUXInst_10_U2  ( .A(AddKey), .B(StateRegOutput[10]), .Z(
        AddKeyMUX_MUXInst_10_n2 ) );
  ORN2 AddKeyMUX_MUXInst_10_U1  ( .A(AddKeyMUX_MUXInst_10_n1 ), .B(
        AddKeyMUX_MUXInst_10_n2 ), .Z(AddKeyMUXOutput[10]) );
  AND2 AddKeyMUX_MUXInst_11_U3  ( .A(Ciphertext[11]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_11_n1 ) );
  ORN2 AddKeyMUX_MUXInst_11_U2  ( .A(AddKey), .B(StateRegOutput[11]), .Z(
        AddKeyMUX_MUXInst_11_n2 ) );
  ORN2 AddKeyMUX_MUXInst_11_U1  ( .A(AddKeyMUX_MUXInst_11_n1 ), .B(
        AddKeyMUX_MUXInst_11_n2 ), .Z(AddKeyMUXOutput[11]) );
  AND2 AddKeyMUX_MUXInst_12_U3  ( .A(Ciphertext[12]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_12_n1 ) );
  ORN2 AddKeyMUX_MUXInst_12_U2  ( .A(AddKey), .B(StateRegOutput[12]), .Z(
        AddKeyMUX_MUXInst_12_n2 ) );
  ORN2 AddKeyMUX_MUXInst_12_U1  ( .A(AddKeyMUX_MUXInst_12_n1 ), .B(
        AddKeyMUX_MUXInst_12_n2 ), .Z(AddKeyMUXOutput[12]) );
  AND2 AddKeyMUX_MUXInst_13_U3  ( .A(Ciphertext[13]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_13_n1 ) );
  ORN2 AddKeyMUX_MUXInst_13_U2  ( .A(AddKey), .B(StateRegOutput[13]), .Z(
        AddKeyMUX_MUXInst_13_n2 ) );
  ORN2 AddKeyMUX_MUXInst_13_U1  ( .A(AddKeyMUX_MUXInst_13_n1 ), .B(
        AddKeyMUX_MUXInst_13_n2 ), .Z(AddKeyMUXOutput[13]) );
  AND2 AddKeyMUX_MUXInst_14_U3  ( .A(Ciphertext[14]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_14_n1 ) );
  ORN2 AddKeyMUX_MUXInst_14_U2  ( .A(AddKey), .B(StateRegOutput[14]), .Z(
        AddKeyMUX_MUXInst_14_n2 ) );
  ORN2 AddKeyMUX_MUXInst_14_U1  ( .A(AddKeyMUX_MUXInst_14_n1 ), .B(
        AddKeyMUX_MUXInst_14_n2 ), .Z(AddKeyMUXOutput[14]) );
  AND2 AddKeyMUX_MUXInst_15_U3  ( .A(Ciphertext[15]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_15_n1 ) );
  ORN2 AddKeyMUX_MUXInst_15_U2  ( .A(AddKey), .B(StateRegOutput[15]), .Z(
        AddKeyMUX_MUXInst_15_n2 ) );
  ORN2 AddKeyMUX_MUXInst_15_U1  ( .A(AddKeyMUX_MUXInst_15_n1 ), .B(
        AddKeyMUX_MUXInst_15_n2 ), .Z(AddKeyMUXOutput[15]) );
  AND2 AddKeyMUX_MUXInst_16_U3  ( .A(Ciphertext[16]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_16_n1 ) );
  ORN2 AddKeyMUX_MUXInst_16_U2  ( .A(AddKey), .B(StateRegOutput[16]), .Z(
        AddKeyMUX_MUXInst_16_n2 ) );
  ORN2 AddKeyMUX_MUXInst_16_U1  ( .A(AddKeyMUX_MUXInst_16_n1 ), .B(
        AddKeyMUX_MUXInst_16_n2 ), .Z(AddKeyMUXOutput[16]) );
  AND2 AddKeyMUX_MUXInst_17_U3  ( .A(Ciphertext[17]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_17_n1 ) );
  ORN2 AddKeyMUX_MUXInst_17_U2  ( .A(AddKey), .B(StateRegOutput[17]), .Z(
        AddKeyMUX_MUXInst_17_n2 ) );
  ORN2 AddKeyMUX_MUXInst_17_U1  ( .A(AddKeyMUX_MUXInst_17_n1 ), .B(
        AddKeyMUX_MUXInst_17_n2 ), .Z(AddKeyMUXOutput[17]) );
  AND2 AddKeyMUX_MUXInst_18_U3  ( .A(Ciphertext[18]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_18_n1 ) );
  ORN2 AddKeyMUX_MUXInst_18_U2  ( .A(AddKey), .B(StateRegOutput[18]), .Z(
        AddKeyMUX_MUXInst_18_n2 ) );
  ORN2 AddKeyMUX_MUXInst_18_U1  ( .A(AddKeyMUX_MUXInst_18_n1 ), .B(
        AddKeyMUX_MUXInst_18_n2 ), .Z(AddKeyMUXOutput[18]) );
  AND2 AddKeyMUX_MUXInst_19_U3  ( .A(Ciphertext[19]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_19_n1 ) );
  ORN2 AddKeyMUX_MUXInst_19_U2  ( .A(AddKey), .B(StateRegOutput[19]), .Z(
        AddKeyMUX_MUXInst_19_n2 ) );
  ORN2 AddKeyMUX_MUXInst_19_U1  ( .A(AddKeyMUX_MUXInst_19_n1 ), .B(
        AddKeyMUX_MUXInst_19_n2 ), .Z(AddKeyMUXOutput[19]) );
  AND2 AddKeyMUX_MUXInst_20_U3  ( .A(Ciphertext[20]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_20_n1 ) );
  ORN2 AddKeyMUX_MUXInst_20_U2  ( .A(AddKey), .B(StateRegOutput[20]), .Z(
        AddKeyMUX_MUXInst_20_n2 ) );
  ORN2 AddKeyMUX_MUXInst_20_U1  ( .A(AddKeyMUX_MUXInst_20_n1 ), .B(
        AddKeyMUX_MUXInst_20_n2 ), .Z(AddKeyMUXOutput[20]) );
  AND2 AddKeyMUX_MUXInst_21_U3  ( .A(Ciphertext[21]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_21_n1 ) );
  ORN2 AddKeyMUX_MUXInst_21_U2  ( .A(AddKey), .B(StateRegOutput[21]), .Z(
        AddKeyMUX_MUXInst_21_n2 ) );
  ORN2 AddKeyMUX_MUXInst_21_U1  ( .A(AddKeyMUX_MUXInst_21_n1 ), .B(
        AddKeyMUX_MUXInst_21_n2 ), .Z(AddKeyMUXOutput[21]) );
  AND2 AddKeyMUX_MUXInst_22_U3  ( .A(Ciphertext[22]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_22_n1 ) );
  ORN2 AddKeyMUX_MUXInst_22_U2  ( .A(AddKey), .B(StateRegOutput[22]), .Z(
        AddKeyMUX_MUXInst_22_n2 ) );
  ORN2 AddKeyMUX_MUXInst_22_U1  ( .A(AddKeyMUX_MUXInst_22_n1 ), .B(
        AddKeyMUX_MUXInst_22_n2 ), .Z(AddKeyMUXOutput[22]) );
  AND2 AddKeyMUX_MUXInst_23_U3  ( .A(Ciphertext[23]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_23_n1 ) );
  ORN2 AddKeyMUX_MUXInst_23_U2  ( .A(AddKey), .B(StateRegOutput[23]), .Z(
        AddKeyMUX_MUXInst_23_n2 ) );
  ORN2 AddKeyMUX_MUXInst_23_U1  ( .A(AddKeyMUX_MUXInst_23_n1 ), .B(
        AddKeyMUX_MUXInst_23_n2 ), .Z(AddKeyMUXOutput[23]) );
  AND2 AddKeyMUX_MUXInst_24_U3  ( .A(Ciphertext[24]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_24_n1 ) );
  ORN2 AddKeyMUX_MUXInst_24_U2  ( .A(AddKey), .B(StateRegOutput[24]), .Z(
        AddKeyMUX_MUXInst_24_n2 ) );
  ORN2 AddKeyMUX_MUXInst_24_U1  ( .A(AddKeyMUX_MUXInst_24_n1 ), .B(
        AddKeyMUX_MUXInst_24_n2 ), .Z(AddKeyMUXOutput[24]) );
  AND2 AddKeyMUX_MUXInst_25_U3  ( .A(Ciphertext[25]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_25_n1 ) );
  ORN2 AddKeyMUX_MUXInst_25_U2  ( .A(AddKey), .B(StateRegOutput[25]), .Z(
        AddKeyMUX_MUXInst_25_n2 ) );
  ORN2 AddKeyMUX_MUXInst_25_U1  ( .A(AddKeyMUX_MUXInst_25_n1 ), .B(
        AddKeyMUX_MUXInst_25_n2 ), .Z(AddKeyMUXOutput[25]) );
  AND2 AddKeyMUX_MUXInst_26_U3  ( .A(Ciphertext[26]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_26_n1 ) );
  ORN2 AddKeyMUX_MUXInst_26_U2  ( .A(AddKey), .B(StateRegOutput[26]), .Z(
        AddKeyMUX_MUXInst_26_n2 ) );
  ORN2 AddKeyMUX_MUXInst_26_U1  ( .A(AddKeyMUX_MUXInst_26_n1 ), .B(
        AddKeyMUX_MUXInst_26_n2 ), .Z(AddKeyMUXOutput[26]) );
  AND2 AddKeyMUX_MUXInst_27_U3  ( .A(Ciphertext[27]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_27_n1 ) );
  ORN2 AddKeyMUX_MUXInst_27_U2  ( .A(AddKey), .B(StateRegOutput[27]), .Z(
        AddKeyMUX_MUXInst_27_n2 ) );
  ORN2 AddKeyMUX_MUXInst_27_U1  ( .A(AddKeyMUX_MUXInst_27_n1 ), .B(
        AddKeyMUX_MUXInst_27_n2 ), .Z(AddKeyMUXOutput[27]) );
  AND2 AddKeyMUX_MUXInst_28_U3  ( .A(Ciphertext[28]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_28_n1 ) );
  ORN2 AddKeyMUX_MUXInst_28_U2  ( .A(AddKey), .B(StateRegOutput[28]), .Z(
        AddKeyMUX_MUXInst_28_n2 ) );
  ORN2 AddKeyMUX_MUXInst_28_U1  ( .A(AddKeyMUX_MUXInst_28_n1 ), .B(
        AddKeyMUX_MUXInst_28_n2 ), .Z(AddKeyMUXOutput[28]) );
  AND2 AddKeyMUX_MUXInst_29_U3  ( .A(Ciphertext[29]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_29_n1 ) );
  ORN2 AddKeyMUX_MUXInst_29_U2  ( .A(AddKey), .B(StateRegOutput[29]), .Z(
        AddKeyMUX_MUXInst_29_n2 ) );
  ORN2 AddKeyMUX_MUXInst_29_U1  ( .A(AddKeyMUX_MUXInst_29_n1 ), .B(
        AddKeyMUX_MUXInst_29_n2 ), .Z(AddKeyMUXOutput[29]) );
  AND2 AddKeyMUX_MUXInst_30_U3  ( .A(Ciphertext[30]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_30_n1 ) );
  ORN2 AddKeyMUX_MUXInst_30_U2  ( .A(AddKey), .B(StateRegOutput[30]), .Z(
        AddKeyMUX_MUXInst_30_n2 ) );
  ORN2 AddKeyMUX_MUXInst_30_U1  ( .A(AddKeyMUX_MUXInst_30_n1 ), .B(
        AddKeyMUX_MUXInst_30_n2 ), .Z(AddKeyMUXOutput[30]) );
  AND2 AddKeyMUX_MUXInst_31_U3  ( .A(Ciphertext[31]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_31_n1 ) );
  ORN2 AddKeyMUX_MUXInst_31_U2  ( .A(AddKey), .B(StateRegOutput[31]), .Z(
        AddKeyMUX_MUXInst_31_n2 ) );
  ORN2 AddKeyMUX_MUXInst_31_U1  ( .A(AddKeyMUX_MUXInst_31_n1 ), .B(
        AddKeyMUX_MUXInst_31_n2 ), .Z(AddKeyMUXOutput[31]) );
  AND2 AddKeyMUX_MUXInst_32_U3  ( .A(Ciphertext[32]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_32_n1 ) );
  ORN2 AddKeyMUX_MUXInst_32_U2  ( .A(AddKey), .B(StateRegOutput[32]), .Z(
        AddKeyMUX_MUXInst_32_n2 ) );
  ORN2 AddKeyMUX_MUXInst_32_U1  ( .A(AddKeyMUX_MUXInst_32_n1 ), .B(
        AddKeyMUX_MUXInst_32_n2 ), .Z(AddKeyMUXOutput[32]) );
  AND2 AddKeyMUX_MUXInst_33_U3  ( .A(Ciphertext[33]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_33_n1 ) );
  ORN2 AddKeyMUX_MUXInst_33_U2  ( .A(AddKey), .B(StateRegOutput[33]), .Z(
        AddKeyMUX_MUXInst_33_n2 ) );
  ORN2 AddKeyMUX_MUXInst_33_U1  ( .A(AddKeyMUX_MUXInst_33_n1 ), .B(
        AddKeyMUX_MUXInst_33_n2 ), .Z(AddKeyMUXOutput[33]) );
  AND2 AddKeyMUX_MUXInst_34_U3  ( .A(Ciphertext[34]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_34_n1 ) );
  ORN2 AddKeyMUX_MUXInst_34_U2  ( .A(AddKey), .B(StateRegOutput[34]), .Z(
        AddKeyMUX_MUXInst_34_n2 ) );
  ORN2 AddKeyMUX_MUXInst_34_U1  ( .A(AddKeyMUX_MUXInst_34_n1 ), .B(
        AddKeyMUX_MUXInst_34_n2 ), .Z(AddKeyMUXOutput[34]) );
  AND2 AddKeyMUX_MUXInst_35_U3  ( .A(Ciphertext[35]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_35_n1 ) );
  ORN2 AddKeyMUX_MUXInst_35_U2  ( .A(AddKey), .B(StateRegOutput[35]), .Z(
        AddKeyMUX_MUXInst_35_n2 ) );
  ORN2 AddKeyMUX_MUXInst_35_U1  ( .A(AddKeyMUX_MUXInst_35_n1 ), .B(
        AddKeyMUX_MUXInst_35_n2 ), .Z(AddKeyMUXOutput[35]) );
  AND2 AddKeyMUX_MUXInst_36_U3  ( .A(Ciphertext[36]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_36_n1 ) );
  ORN2 AddKeyMUX_MUXInst_36_U2  ( .A(AddKey), .B(StateRegOutput[36]), .Z(
        AddKeyMUX_MUXInst_36_n2 ) );
  ORN2 AddKeyMUX_MUXInst_36_U1  ( .A(AddKeyMUX_MUXInst_36_n1 ), .B(
        AddKeyMUX_MUXInst_36_n2 ), .Z(AddKeyMUXOutput[36]) );
  AND2 AddKeyMUX_MUXInst_37_U3  ( .A(Ciphertext[37]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_37_n1 ) );
  ORN2 AddKeyMUX_MUXInst_37_U2  ( .A(AddKey), .B(StateRegOutput[37]), .Z(
        AddKeyMUX_MUXInst_37_n2 ) );
  ORN2 AddKeyMUX_MUXInst_37_U1  ( .A(AddKeyMUX_MUXInst_37_n1 ), .B(
        AddKeyMUX_MUXInst_37_n2 ), .Z(AddKeyMUXOutput[37]) );
  AND2 AddKeyMUX_MUXInst_38_U3  ( .A(Ciphertext[38]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_38_n1 ) );
  ORN2 AddKeyMUX_MUXInst_38_U2  ( .A(AddKey), .B(StateRegOutput[38]), .Z(
        AddKeyMUX_MUXInst_38_n2 ) );
  ORN2 AddKeyMUX_MUXInst_38_U1  ( .A(AddKeyMUX_MUXInst_38_n1 ), .B(
        AddKeyMUX_MUXInst_38_n2 ), .Z(AddKeyMUXOutput[38]) );
  AND2 AddKeyMUX_MUXInst_39_U3  ( .A(Ciphertext[39]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_39_n1 ) );
  ORN2 AddKeyMUX_MUXInst_39_U2  ( .A(AddKey), .B(StateRegOutput[39]), .Z(
        AddKeyMUX_MUXInst_39_n2 ) );
  ORN2 AddKeyMUX_MUXInst_39_U1  ( .A(AddKeyMUX_MUXInst_39_n1 ), .B(
        AddKeyMUX_MUXInst_39_n2 ), .Z(AddKeyMUXOutput[39]) );
  AND2 AddKeyMUX_MUXInst_40_U3  ( .A(Ciphertext[40]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_40_n1 ) );
  ORN2 AddKeyMUX_MUXInst_40_U2  ( .A(AddKey), .B(StateRegOutput[40]), .Z(
        AddKeyMUX_MUXInst_40_n2 ) );
  ORN2 AddKeyMUX_MUXInst_40_U1  ( .A(AddKeyMUX_MUXInst_40_n1 ), .B(
        AddKeyMUX_MUXInst_40_n2 ), .Z(AddKeyMUXOutput[40]) );
  AND2 AddKeyMUX_MUXInst_41_U3  ( .A(Ciphertext[41]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_41_n1 ) );
  ORN2 AddKeyMUX_MUXInst_41_U2  ( .A(AddKey), .B(StateRegOutput[41]), .Z(
        AddKeyMUX_MUXInst_41_n2 ) );
  ORN2 AddKeyMUX_MUXInst_41_U1  ( .A(AddKeyMUX_MUXInst_41_n1 ), .B(
        AddKeyMUX_MUXInst_41_n2 ), .Z(AddKeyMUXOutput[41]) );
  AND2 AddKeyMUX_MUXInst_42_U3  ( .A(Ciphertext[42]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_42_n1 ) );
  ORN2 AddKeyMUX_MUXInst_42_U2  ( .A(AddKey), .B(StateRegOutput[42]), .Z(
        AddKeyMUX_MUXInst_42_n2 ) );
  ORN2 AddKeyMUX_MUXInst_42_U1  ( .A(AddKeyMUX_MUXInst_42_n1 ), .B(
        AddKeyMUX_MUXInst_42_n2 ), .Z(AddKeyMUXOutput[42]) );
  AND2 AddKeyMUX_MUXInst_43_U3  ( .A(Ciphertext[43]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_43_n1 ) );
  ORN2 AddKeyMUX_MUXInst_43_U2  ( .A(AddKey), .B(StateRegOutput[43]), .Z(
        AddKeyMUX_MUXInst_43_n2 ) );
  ORN2 AddKeyMUX_MUXInst_43_U1  ( .A(AddKeyMUX_MUXInst_43_n1 ), .B(
        AddKeyMUX_MUXInst_43_n2 ), .Z(AddKeyMUXOutput[43]) );
  AND2 AddKeyMUX_MUXInst_44_U3  ( .A(Ciphertext[44]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_44_n1 ) );
  ORN2 AddKeyMUX_MUXInst_44_U2  ( .A(AddKey), .B(StateRegOutput[44]), .Z(
        AddKeyMUX_MUXInst_44_n2 ) );
  ORN2 AddKeyMUX_MUXInst_44_U1  ( .A(AddKeyMUX_MUXInst_44_n1 ), .B(
        AddKeyMUX_MUXInst_44_n2 ), .Z(AddKeyMUXOutput[44]) );
  AND2 AddKeyMUX_MUXInst_45_U3  ( .A(Ciphertext[45]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_45_n1 ) );
  ORN2 AddKeyMUX_MUXInst_45_U2  ( .A(AddKey), .B(StateRegOutput[45]), .Z(
        AddKeyMUX_MUXInst_45_n2 ) );
  ORN2 AddKeyMUX_MUXInst_45_U1  ( .A(AddKeyMUX_MUXInst_45_n1 ), .B(
        AddKeyMUX_MUXInst_45_n2 ), .Z(AddKeyMUXOutput[45]) );
  AND2 AddKeyMUX_MUXInst_46_U3  ( .A(Ciphertext[46]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_46_n1 ) );
  ORN2 AddKeyMUX_MUXInst_46_U2  ( .A(AddKey), .B(StateRegOutput[46]), .Z(
        AddKeyMUX_MUXInst_46_n2 ) );
  ORN2 AddKeyMUX_MUXInst_46_U1  ( .A(AddKeyMUX_MUXInst_46_n1 ), .B(
        AddKeyMUX_MUXInst_46_n2 ), .Z(AddKeyMUXOutput[46]) );
  AND2 AddKeyMUX_MUXInst_47_U3  ( .A(Ciphertext[47]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_47_n1 ) );
  ORN2 AddKeyMUX_MUXInst_47_U2  ( .A(AddKey), .B(StateRegOutput[47]), .Z(
        AddKeyMUX_MUXInst_47_n2 ) );
  ORN2 AddKeyMUX_MUXInst_47_U1  ( .A(AddKeyMUX_MUXInst_47_n1 ), .B(
        AddKeyMUX_MUXInst_47_n2 ), .Z(AddKeyMUXOutput[47]) );
  AND2 AddKeyMUX_MUXInst_48_U3  ( .A(Ciphertext[48]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_48_n1 ) );
  ORN2 AddKeyMUX_MUXInst_48_U2  ( .A(AddKey), .B(StateRegOutput[48]), .Z(
        AddKeyMUX_MUXInst_48_n2 ) );
  ORN2 AddKeyMUX_MUXInst_48_U1  ( .A(AddKeyMUX_MUXInst_48_n1 ), .B(
        AddKeyMUX_MUXInst_48_n2 ), .Z(AddKeyMUXOutput[48]) );
  AND2 AddKeyMUX_MUXInst_49_U3  ( .A(Ciphertext[49]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_49_n1 ) );
  ORN2 AddKeyMUX_MUXInst_49_U2  ( .A(AddKey), .B(StateRegOutput[49]), .Z(
        AddKeyMUX_MUXInst_49_n2 ) );
  ORN2 AddKeyMUX_MUXInst_49_U1  ( .A(AddKeyMUX_MUXInst_49_n1 ), .B(
        AddKeyMUX_MUXInst_49_n2 ), .Z(AddKeyMUXOutput[49]) );
  AND2 AddKeyMUX_MUXInst_50_U3  ( .A(Ciphertext[50]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_50_n1 ) );
  ORN2 AddKeyMUX_MUXInst_50_U2  ( .A(AddKey), .B(StateRegOutput[50]), .Z(
        AddKeyMUX_MUXInst_50_n2 ) );
  ORN2 AddKeyMUX_MUXInst_50_U1  ( .A(AddKeyMUX_MUXInst_50_n1 ), .B(
        AddKeyMUX_MUXInst_50_n2 ), .Z(AddKeyMUXOutput[50]) );
  AND2 AddKeyMUX_MUXInst_51_U3  ( .A(Ciphertext[51]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_51_n1 ) );
  ORN2 AddKeyMUX_MUXInst_51_U2  ( .A(AddKey), .B(StateRegOutput[51]), .Z(
        AddKeyMUX_MUXInst_51_n2 ) );
  ORN2 AddKeyMUX_MUXInst_51_U1  ( .A(AddKeyMUX_MUXInst_51_n1 ), .B(
        AddKeyMUX_MUXInst_51_n2 ), .Z(AddKeyMUXOutput[51]) );
  AND2 AddKeyMUX_MUXInst_52_U3  ( .A(Ciphertext[52]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_52_n1 ) );
  ORN2 AddKeyMUX_MUXInst_52_U2  ( .A(AddKey), .B(StateRegOutput[52]), .Z(
        AddKeyMUX_MUXInst_52_n2 ) );
  ORN2 AddKeyMUX_MUXInst_52_U1  ( .A(AddKeyMUX_MUXInst_52_n1 ), .B(
        AddKeyMUX_MUXInst_52_n2 ), .Z(AddKeyMUXOutput[52]) );
  AND2 AddKeyMUX_MUXInst_53_U3  ( .A(Ciphertext[53]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_53_n1 ) );
  ORN2 AddKeyMUX_MUXInst_53_U2  ( .A(AddKey), .B(StateRegOutput[53]), .Z(
        AddKeyMUX_MUXInst_53_n2 ) );
  ORN2 AddKeyMUX_MUXInst_53_U1  ( .A(AddKeyMUX_MUXInst_53_n1 ), .B(
        AddKeyMUX_MUXInst_53_n2 ), .Z(AddKeyMUXOutput[53]) );
  AND2 AddKeyMUX_MUXInst_54_U3  ( .A(Ciphertext[54]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_54_n1 ) );
  ORN2 AddKeyMUX_MUXInst_54_U2  ( .A(AddKey), .B(StateRegOutput[54]), .Z(
        AddKeyMUX_MUXInst_54_n2 ) );
  ORN2 AddKeyMUX_MUXInst_54_U1  ( .A(AddKeyMUX_MUXInst_54_n1 ), .B(
        AddKeyMUX_MUXInst_54_n2 ), .Z(AddKeyMUXOutput[54]) );
  AND2 AddKeyMUX_MUXInst_55_U3  ( .A(Ciphertext[55]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_55_n1 ) );
  ORN2 AddKeyMUX_MUXInst_55_U2  ( .A(AddKey), .B(StateRegOutput[55]), .Z(
        AddKeyMUX_MUXInst_55_n2 ) );
  ORN2 AddKeyMUX_MUXInst_55_U1  ( .A(AddKeyMUX_MUXInst_55_n1 ), .B(
        AddKeyMUX_MUXInst_55_n2 ), .Z(AddKeyMUXOutput[55]) );
  AND2 AddKeyMUX_MUXInst_56_U3  ( .A(Ciphertext[56]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_56_n1 ) );
  ORN2 AddKeyMUX_MUXInst_56_U2  ( .A(AddKey), .B(StateRegOutput[56]), .Z(
        AddKeyMUX_MUXInst_56_n2 ) );
  ORN2 AddKeyMUX_MUXInst_56_U1  ( .A(AddKeyMUX_MUXInst_56_n1 ), .B(
        AddKeyMUX_MUXInst_56_n2 ), .Z(AddKeyMUXOutput[56]) );
  AND2 AddKeyMUX_MUXInst_57_U3  ( .A(Ciphertext[57]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_57_n1 ) );
  ORN2 AddKeyMUX_MUXInst_57_U2  ( .A(AddKey), .B(StateRegOutput[57]), .Z(
        AddKeyMUX_MUXInst_57_n2 ) );
  ORN2 AddKeyMUX_MUXInst_57_U1  ( .A(AddKeyMUX_MUXInst_57_n1 ), .B(
        AddKeyMUX_MUXInst_57_n2 ), .Z(AddKeyMUXOutput[57]) );
  AND2 AddKeyMUX_MUXInst_58_U3  ( .A(Ciphertext[58]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_58_n1 ) );
  ORN2 AddKeyMUX_MUXInst_58_U2  ( .A(AddKey), .B(StateRegOutput[58]), .Z(
        AddKeyMUX_MUXInst_58_n2 ) );
  ORN2 AddKeyMUX_MUXInst_58_U1  ( .A(AddKeyMUX_MUXInst_58_n1 ), .B(
        AddKeyMUX_MUXInst_58_n2 ), .Z(AddKeyMUXOutput[58]) );
  AND2 AddKeyMUX_MUXInst_59_U3  ( .A(Ciphertext[59]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_59_n1 ) );
  ORN2 AddKeyMUX_MUXInst_59_U2  ( .A(AddKey), .B(StateRegOutput[59]), .Z(
        AddKeyMUX_MUXInst_59_n2 ) );
  ORN2 AddKeyMUX_MUXInst_59_U1  ( .A(AddKeyMUX_MUXInst_59_n1 ), .B(
        AddKeyMUX_MUXInst_59_n2 ), .Z(AddKeyMUXOutput[59]) );
  AND2 AddKeyMUX_MUXInst_60_U3  ( .A(Ciphertext[60]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_60_n1 ) );
  ORN2 AddKeyMUX_MUXInst_60_U2  ( .A(AddKey), .B(StateRegOutput[60]), .Z(
        AddKeyMUX_MUXInst_60_n2 ) );
  ORN2 AddKeyMUX_MUXInst_60_U1  ( .A(AddKeyMUX_MUXInst_60_n1 ), .B(
        AddKeyMUX_MUXInst_60_n2 ), .Z(AddKeyMUXOutput[60]) );
  AND2 AddKeyMUX_MUXInst_61_U3  ( .A(Ciphertext[61]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_61_n1 ) );
  ORN2 AddKeyMUX_MUXInst_61_U2  ( .A(AddKey), .B(StateRegOutput[61]), .Z(
        AddKeyMUX_MUXInst_61_n2 ) );
  ORN2 AddKeyMUX_MUXInst_61_U1  ( .A(AddKeyMUX_MUXInst_61_n1 ), .B(
        AddKeyMUX_MUXInst_61_n2 ), .Z(AddKeyMUXOutput[61]) );
  AND2 AddKeyMUX_MUXInst_62_U3  ( .A(Ciphertext[62]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_62_n1 ) );
  ORN2 AddKeyMUX_MUXInst_62_U2  ( .A(AddKey), .B(StateRegOutput[62]), .Z(
        AddKeyMUX_MUXInst_62_n2 ) );
  ORN2 AddKeyMUX_MUXInst_62_U1  ( .A(AddKeyMUX_MUXInst_62_n1 ), .B(
        AddKeyMUX_MUXInst_62_n2 ), .Z(AddKeyMUXOutput[62]) );
  AND2 AddKeyMUX_MUXInst_63_U3  ( .A(Ciphertext[63]), .B(AddKey), .Z(
        AddKeyMUX_MUXInst_63_n1 ) );
  ORN2 AddKeyMUX_MUXInst_63_U2  ( .A(AddKey), .B(StateRegOutput[63]), .Z(
        AddKeyMUX_MUXInst_63_n2 ) );
  ORN2 AddKeyMUX_MUXInst_63_U1  ( .A(AddKeyMUX_MUXInst_63_n1 ), .B(
        AddKeyMUX_MUXInst_63_n2 ), .Z(AddKeyMUXOutput[63]) );
  XOR2 AddConstXOR_XORInst_XORInst_0_0_U2  ( .A(FSMUpdate[1]), .B(
        AddKeyMUXOutput[8]), .Z(AddConstXOR_XORInst_XORInst_0_0_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_0_0_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_0_0_n1 ), .Z(AddConstOutput[0]) );
  XOR2 AddConstXOR_XORInst_XORInst_0_1_U2  ( .A(FSM[1]), .B(
        AddKeyMUXOutput[9]), .Z(AddConstXOR_XORInst_XORInst_0_1_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_0_1_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_0_1_n1 ), .Z(AddConstOutput[1]) );
  XOR2 AddConstXOR_XORInst_XORInst_0_2_U2  ( .A(FSMUpdate[3]), .B(
        AddKeyMUXOutput[10]), .Z(AddConstXOR_XORInst_XORInst_0_2_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_0_2_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_0_2_n1 ), .Z(AddConstOutput[2]) );
  XOR2 AddConstXOR_XORInst_XORInst_0_3_U2  ( .A(1'b0), .B(AddKeyMUXOutput[11]), .Z(AddConstXOR_XORInst_XORInst_0_3_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_0_3_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_0_3_n1 ), .Z(AddConstOutput[3]) );
  XOR2 AddConstXOR_XORInst_XORInst_1_0_U2  ( .A(1'b1), .B(AddKeyMUXOutput[12]), .Z(AddConstXOR_XORInst_XORInst_1_0_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_1_0_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_1_0_n1 ), .Z(AddConstOutput[4]) );
  XOR2 AddConstXOR_XORInst_XORInst_1_1_U2  ( .A(1'b1), .B(AddKeyMUXOutput[13]), .Z(AddConstXOR_XORInst_XORInst_1_1_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_1_1_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_1_1_n1 ), .Z(AddConstOutput[5]) );
  XOR2 AddConstXOR_XORInst_XORInst_1_2_U2  ( .A(1'b0), .B(AddKeyMUXOutput[14]), .Z(AddConstXOR_XORInst_XORInst_1_2_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_1_2_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_1_2_n1 ), .Z(AddConstOutput[6]) );
  XOR2 AddConstXOR_XORInst_XORInst_1_3_U2  ( .A(1'b0), .B(AddKeyMUXOutput[15]), .Z(AddConstXOR_XORInst_XORInst_1_3_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_1_3_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_1_3_n1 ), .Z(AddConstOutput[7]) );
  XOR2 AddConstXOR_XORInst_XORInst_2_0_U2  ( .A(FSMUpdate[4]), .B(
        AddKeyMUXOutput[24]), .Z(AddConstXOR_XORInst_XORInst_2_0_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_2_0_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_2_0_n1 ), .Z(AddConstOutput[8]) );
  XOR2 AddConstXOR_XORInst_XORInst_2_1_U2  ( .A(FSM[4]), .B(
        AddKeyMUXOutput[25]), .Z(AddConstXOR_XORInst_XORInst_2_1_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_2_1_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_2_1_n1 ), .Z(AddConstOutput[9]) );
  XOR2 AddConstXOR_XORInst_XORInst_2_2_U2  ( .A(FSM[5]), .B(
        AddKeyMUXOutput[26]), .Z(AddConstXOR_XORInst_XORInst_2_2_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_2_2_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_2_2_n1 ), .Z(AddConstOutput[10]) );
  XOR2 AddConstXOR_XORInst_XORInst_2_3_U2  ( .A(1'b0), .B(AddKeyMUXOutput[27]), .Z(AddConstXOR_XORInst_XORInst_2_3_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_2_3_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_2_3_n1 ), .Z(AddConstOutput[11]) );
  XOR2 AddConstXOR_XORInst_XORInst_3_0_U2  ( .A(1'b0), .B(AddKeyMUXOutput[28]), .Z(AddConstXOR_XORInst_XORInst_3_0_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_3_0_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_3_0_n1 ), .Z(AddConstOutput[12]) );
  XOR2 AddConstXOR_XORInst_XORInst_3_1_U2  ( .A(1'b1), .B(AddKeyMUXOutput[29]), .Z(AddConstXOR_XORInst_XORInst_3_1_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_3_1_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_3_1_n1 ), .Z(AddConstOutput[13]) );
  XOR2 AddConstXOR_XORInst_XORInst_3_2_U2  ( .A(1'b0), .B(AddKeyMUXOutput[30]), .Z(AddConstXOR_XORInst_XORInst_3_2_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_3_2_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_3_2_n1 ), .Z(AddConstOutput[14]) );
  XOR2 AddConstXOR_XORInst_XORInst_3_3_U2  ( .A(1'b0), .B(AddKeyMUXOutput[31]), .Z(AddConstXOR_XORInst_XORInst_3_3_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_3_3_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_3_3_n1 ), .Z(AddConstOutput[15]) );
  XOR2 AddConstXOR_XORInst_XORInst_4_0_U2  ( .A(FSMUpdate[1]), .B(
        AddKeyMUXOutput[40]), .Z(AddConstXOR_XORInst_XORInst_4_0_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_4_0_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_4_0_n1 ), .Z(AddConstOutput[16]) );
  XOR2 AddConstXOR_XORInst_XORInst_4_1_U2  ( .A(FSM[1]), .B(
        AddKeyMUXOutput[41]), .Z(AddConstXOR_XORInst_XORInst_4_1_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_4_1_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_4_1_n1 ), .Z(AddConstOutput[17]) );
  XOR2 AddConstXOR_XORInst_XORInst_4_2_U2  ( .A(FSMUpdate[3]), .B(
        AddKeyMUXOutput[42]), .Z(AddConstXOR_XORInst_XORInst_4_2_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_4_2_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_4_2_n1 ), .Z(AddConstOutput[18]) );
  XOR2 AddConstXOR_XORInst_XORInst_4_3_U2  ( .A(1'b0), .B(AddKeyMUXOutput[43]), .Z(AddConstXOR_XORInst_XORInst_4_3_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_4_3_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_4_3_n1 ), .Z(AddConstOutput[19]) );
  XOR2 AddConstXOR_XORInst_XORInst_5_0_U2  ( .A(1'b1), .B(AddKeyMUXOutput[44]), .Z(AddConstXOR_XORInst_XORInst_5_0_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_5_0_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_5_0_n1 ), .Z(AddConstOutput[20]) );
  XOR2 AddConstXOR_XORInst_XORInst_5_1_U2  ( .A(1'b0), .B(AddKeyMUXOutput[45]), .Z(AddConstXOR_XORInst_XORInst_5_1_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_5_1_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_5_1_n1 ), .Z(AddConstOutput[21]) );
  XOR2 AddConstXOR_XORInst_XORInst_5_2_U2  ( .A(1'b1), .B(AddKeyMUXOutput[46]), .Z(AddConstXOR_XORInst_XORInst_5_2_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_5_2_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_5_2_n1 ), .Z(AddConstOutput[22]) );
  XOR2 AddConstXOR_XORInst_XORInst_5_3_U2  ( .A(1'b0), .B(AddKeyMUXOutput[47]), .Z(AddConstXOR_XORInst_XORInst_5_3_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_5_3_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_5_3_n1 ), .Z(AddConstOutput[23]) );
  XOR2 AddConstXOR_XORInst_XORInst_6_0_U2  ( .A(FSMUpdate[4]), .B(
        AddKeyMUXOutput[56]), .Z(AddConstXOR_XORInst_XORInst_6_0_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_6_0_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_6_0_n1 ), .Z(AddConstOutput[24]) );
  XOR2 AddConstXOR_XORInst_XORInst_6_1_U2  ( .A(FSM[4]), .B(
        AddKeyMUXOutput[57]), .Z(AddConstXOR_XORInst_XORInst_6_1_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_6_1_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_6_1_n1 ), .Z(AddConstOutput[25]) );
  XOR2 AddConstXOR_XORInst_XORInst_6_2_U2  ( .A(FSM[5]), .B(
        AddKeyMUXOutput[58]), .Z(AddConstXOR_XORInst_XORInst_6_2_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_6_2_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_6_2_n1 ), .Z(AddConstOutput[26]) );
  XOR2 AddConstXOR_XORInst_XORInst_6_3_U2  ( .A(1'b0), .B(AddKeyMUXOutput[59]), .Z(AddConstXOR_XORInst_XORInst_6_3_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_6_3_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_6_3_n1 ), .Z(AddConstOutput[27]) );
  XOR2 AddConstXOR_XORInst_XORInst_7_0_U2  ( .A(1'b0), .B(AddKeyMUXOutput[60]), .Z(AddConstXOR_XORInst_XORInst_7_0_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_7_0_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_7_0_n1 ), .Z(AddConstOutput[28]) );
  XOR2 AddConstXOR_XORInst_XORInst_7_1_U2  ( .A(1'b0), .B(AddKeyMUXOutput[61]), .Z(AddConstXOR_XORInst_XORInst_7_1_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_7_1_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_7_1_n1 ), .Z(AddConstOutput[29]) );
  XOR2 AddConstXOR_XORInst_XORInst_7_2_U2  ( .A(1'b1), .B(AddKeyMUXOutput[62]), .Z(AddConstXOR_XORInst_XORInst_7_2_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_7_2_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_7_2_n1 ), .Z(AddConstOutput[30]) );
  XOR2 AddConstXOR_XORInst_XORInst_7_3_U2  ( .A(1'b0), .B(AddKeyMUXOutput[63]), .Z(AddConstXOR_XORInst_XORInst_7_3_n1 ) );
  XOR2 AddConstXOR_XORInst_XORInst_7_3_U1  ( .A(1'b0), .B(
        AddConstXOR_XORInst_XORInst_7_3_n1 ), .Z(AddConstOutput[31]) );
  OR2 SubCellInst_LFInst_0_LFInst_3_U9  ( .A(AddKeyMUXOutput[1]), .B(
        AddKeyMUXOutput[0]), .Z(SubCellInst_LFInst_0_LFInst_3_n5 ) );
  AND2 SubCellInst_LFInst_0_LFInst_3_U8  ( .A(AddKeyMUXOutput[3]), .B(
        SubCellInst_LFInst_0_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_0_LFInst_3_n7 ) );
  AND2 SubCellInst_LFInst_0_LFInst_3_U7  ( .A(AddKeyMUXOutput[0]), .B(
        AddKeyMUXOutput[1]), .Z(SubCellInst_LFInst_0_LFInst_3_n8 ) );
  OR2 SubCellInst_LFInst_0_LFInst_3_U6  ( .A(
        SubCellInst_LFInst_0_LFInst_3_n7 ), .B(
        SubCellInst_LFInst_0_LFInst_3_n8 ), .Z(
        SubCellInst_LFInst_0_LFInst_3_n6 ) );
  BIC2 SubCellInst_LFInst_0_LFInst_3_U5  ( .A(
        SubCellInst_LFInst_0_LFInst_3_n6 ), .B(AddKeyMUXOutput[2]), .Z(
        SubCellInst_LFInst_0_LFInst_3_n1 ) );
  AND2 SubCellInst_LFInst_0_LFInst_3_U4  ( .A(AddKeyMUXOutput[2]), .B(
        AddKeyMUXOutput[1]), .Z(SubCellInst_LFInst_0_LFInst_3_n4 ) );
  ORN2 SubCellInst_LFInst_0_LFInst_3_U3  ( .A(
        SubCellInst_LFInst_0_LFInst_3_n4 ), .B(
        SubCellInst_LFInst_0_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_0_LFInst_3_n3 ) );
  ORN2 SubCellInst_LFInst_0_LFInst_3_U2  ( .A(AddKeyMUXOutput[3]), .B(
        SubCellInst_LFInst_0_LFInst_3_n3 ), .Z(
        SubCellInst_LFInst_0_LFInst_3_n2 ) );
  ORN2 SubCellInst_LFInst_0_LFInst_3_U1  ( .A(
        SubCellInst_LFInst_0_LFInst_3_n1 ), .B(
        SubCellInst_LFInst_0_LFInst_3_n2 ), .Z(MCInst1_MC0_v3_2 [2]) );
  BIC2 SubCellInst_LFInst_0_LFInst_2_U11  ( .A(AddKeyMUXOutput[1]), .B(
        AddKeyMUXOutput[0]), .Z(SubCellInst_LFInst_0_LFInst_2_n8 ) );
  ORN2 SubCellInst_LFInst_0_LFInst_2_U10  ( .A(AddKeyMUXOutput[0]), .B(
        AddKeyMUXOutput[3]), .Z(SubCellInst_LFInst_0_LFInst_2_n10 ) );
  ORN2 SubCellInst_LFInst_0_LFInst_2_U9  ( .A(AddKeyMUXOutput[1]), .B(
        SubCellInst_LFInst_0_LFInst_2_n10 ), .Z(
        SubCellInst_LFInst_0_LFInst_2_n9 ) );
  ORN2 SubCellInst_LFInst_0_LFInst_2_U8  ( .A(
        SubCellInst_LFInst_0_LFInst_2_n8 ), .B(
        SubCellInst_LFInst_0_LFInst_2_n9 ), .Z(
        SubCellInst_LFInst_0_LFInst_2_n7 ) );
  BIC2 SubCellInst_LFInst_0_LFInst_2_U7  ( .A(
        SubCellInst_LFInst_0_LFInst_2_n7 ), .B(AddKeyMUXOutput[2]), .Z(
        SubCellInst_LFInst_0_LFInst_2_n1 ) );
  ORN2 SubCellInst_LFInst_0_LFInst_2_U6  ( .A(AddKeyMUXOutput[1]), .B(
        AddKeyMUXOutput[3]), .Z(SubCellInst_LFInst_0_LFInst_2_n4 ) );
  AND2 SubCellInst_LFInst_0_LFInst_2_U5  ( .A(AddKeyMUXOutput[1]), .B(
        AddKeyMUXOutput[0]), .Z(SubCellInst_LFInst_0_LFInst_2_n6 ) );
  ORN2 SubCellInst_LFInst_0_LFInst_2_U4  ( .A(AddKeyMUXOutput[3]), .B(
        SubCellInst_LFInst_0_LFInst_2_n6 ), .Z(
        SubCellInst_LFInst_0_LFInst_2_n5 ) );
  AND2 SubCellInst_LFInst_0_LFInst_2_U3  ( .A(
        SubCellInst_LFInst_0_LFInst_2_n4 ), .B(
        SubCellInst_LFInst_0_LFInst_2_n5 ), .Z(
        SubCellInst_LFInst_0_LFInst_2_n3 ) );
  ORN2 SubCellInst_LFInst_0_LFInst_2_U2  ( .A(
        SubCellInst_LFInst_0_LFInst_2_n3 ), .B(AddKeyMUXOutput[2]), .Z(
        SubCellInst_LFInst_0_LFInst_2_n2 ) );
  ORN2 SubCellInst_LFInst_0_LFInst_2_U1  ( .A(
        SubCellInst_LFInst_0_LFInst_2_n1 ), .B(
        SubCellInst_LFInst_0_LFInst_2_n2 ), .Z(MCInst1_MC0_v3_0 [3]) );
  AND2 SubCellInst_LFInst_0_LFInst_1_U8  ( .A(AddKeyMUXOutput[2]), .B(
        AddKeyMUXOutput[0]), .Z(SubCellInst_LFInst_0_LFInst_1_n4 ) );
  AND2 SubCellInst_LFInst_0_LFInst_1_U7  ( .A(AddKeyMUXOutput[1]), .B(
        AddKeyMUXOutput[0]), .Z(SubCellInst_LFInst_0_LFInst_1_n7 ) );
  OR2 SubCellInst_LFInst_0_LFInst_1_U6  ( .A(AddKeyMUXOutput[2]), .B(
        SubCellInst_LFInst_0_LFInst_1_n7 ), .Z(
        SubCellInst_LFInst_0_LFInst_1_n6 ) );
  ORN2 SubCellInst_LFInst_0_LFInst_1_U5  ( .A(
        SubCellInst_LFInst_0_LFInst_1_n4 ), .B(
        SubCellInst_LFInst_0_LFInst_1_n6 ), .Z(
        SubCellInst_LFInst_0_LFInst_1_n5 ) );
  AND2 SubCellInst_LFInst_0_LFInst_1_U4  ( .A(AddKeyMUXOutput[3]), .B(
        SubCellInst_LFInst_0_LFInst_1_n5 ), .Z(
        SubCellInst_LFInst_0_LFInst_1_n1 ) );
  BIC2 SubCellInst_LFInst_0_LFInst_1_U3  ( .A(AddKeyMUXOutput[1]), .B(
        SubCellInst_LFInst_0_LFInst_1_n4 ), .Z(
        SubCellInst_LFInst_0_LFInst_1_n3 ) );
  ORN2 SubCellInst_LFInst_0_LFInst_1_U2  ( .A(AddKeyMUXOutput[3]), .B(
        SubCellInst_LFInst_0_LFInst_1_n3 ), .Z(
        SubCellInst_LFInst_0_LFInst_1_n2 ) );
  ORN2 SubCellInst_LFInst_0_LFInst_1_U1  ( .A(
        SubCellInst_LFInst_0_LFInst_1_n1 ), .B(
        SubCellInst_LFInst_0_LFInst_1_n2 ), .Z(MCInst1_MC0_v3_0 [2]) );
  BIC2 SubCellInst_LFInst_0_LFInst_0_U3  ( .A(AddKeyMUXOutput[2]), .B(
        AddKeyMUXOutput[1]), .Z(SubCellInst_LFInst_0_LFInst_0_n1 ) );
  XOR2 SubCellInst_LFInst_0_LFInst_0_U2  ( .A(AddKeyMUXOutput[3]), .B(
        AddKeyMUXOutput[0]), .Z(SubCellInst_LFInst_0_LFInst_0_n2 ) );
  XOR2 SubCellInst_LFInst_0_LFInst_0_U1  ( .A(
        SubCellInst_LFInst_0_LFInst_0_n1 ), .B(
        SubCellInst_LFInst_0_LFInst_0_n2 ), .Z(MCInst1_MC0_v3_2 [3]) );
  OR2 SubCellInst_LFInst_1_LFInst_3_U9  ( .A(AddKeyMUXOutput[5]), .B(
        AddKeyMUXOutput[4]), .Z(SubCellInst_LFInst_1_LFInst_3_n5 ) );
  AND2 SubCellInst_LFInst_1_LFInst_3_U8  ( .A(AddKeyMUXOutput[7]), .B(
        SubCellInst_LFInst_1_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_1_LFInst_3_n7 ) );
  AND2 SubCellInst_LFInst_1_LFInst_3_U7  ( .A(AddKeyMUXOutput[4]), .B(
        AddKeyMUXOutput[5]), .Z(SubCellInst_LFInst_1_LFInst_3_n8 ) );
  OR2 SubCellInst_LFInst_1_LFInst_3_U6  ( .A(
        SubCellInst_LFInst_1_LFInst_3_n7 ), .B(
        SubCellInst_LFInst_1_LFInst_3_n8 ), .Z(
        SubCellInst_LFInst_1_LFInst_3_n6 ) );
  BIC2 SubCellInst_LFInst_1_LFInst_3_U5  ( .A(
        SubCellInst_LFInst_1_LFInst_3_n6 ), .B(AddKeyMUXOutput[6]), .Z(
        SubCellInst_LFInst_1_LFInst_3_n1 ) );
  AND2 SubCellInst_LFInst_1_LFInst_3_U4  ( .A(AddKeyMUXOutput[6]), .B(
        AddKeyMUXOutput[5]), .Z(SubCellInst_LFInst_1_LFInst_3_n4 ) );
  ORN2 SubCellInst_LFInst_1_LFInst_3_U3  ( .A(
        SubCellInst_LFInst_1_LFInst_3_n4 ), .B(
        SubCellInst_LFInst_1_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_1_LFInst_3_n3 ) );
  ORN2 SubCellInst_LFInst_1_LFInst_3_U2  ( .A(AddKeyMUXOutput[7]), .B(
        SubCellInst_LFInst_1_LFInst_3_n3 ), .Z(
        SubCellInst_LFInst_1_LFInst_3_n2 ) );
  ORN2 SubCellInst_LFInst_1_LFInst_3_U1  ( .A(
        SubCellInst_LFInst_1_LFInst_3_n1 ), .B(
        SubCellInst_LFInst_1_LFInst_3_n2 ), .Z(MCInst1_MC3_v3_2 [2]) );
  BIC2 SubCellInst_LFInst_1_LFInst_2_U11  ( .A(AddKeyMUXOutput[5]), .B(
        AddKeyMUXOutput[4]), .Z(SubCellInst_LFInst_1_LFInst_2_n8 ) );
  ORN2 SubCellInst_LFInst_1_LFInst_2_U10  ( .A(AddKeyMUXOutput[4]), .B(
        AddKeyMUXOutput[7]), .Z(SubCellInst_LFInst_1_LFInst_2_n10 ) );
  ORN2 SubCellInst_LFInst_1_LFInst_2_U9  ( .A(AddKeyMUXOutput[5]), .B(
        SubCellInst_LFInst_1_LFInst_2_n10 ), .Z(
        SubCellInst_LFInst_1_LFInst_2_n9 ) );
  ORN2 SubCellInst_LFInst_1_LFInst_2_U8  ( .A(
        SubCellInst_LFInst_1_LFInst_2_n8 ), .B(
        SubCellInst_LFInst_1_LFInst_2_n9 ), .Z(
        SubCellInst_LFInst_1_LFInst_2_n7 ) );
  BIC2 SubCellInst_LFInst_1_LFInst_2_U7  ( .A(
        SubCellInst_LFInst_1_LFInst_2_n7 ), .B(AddKeyMUXOutput[6]), .Z(
        SubCellInst_LFInst_1_LFInst_2_n1 ) );
  ORN2 SubCellInst_LFInst_1_LFInst_2_U6  ( .A(AddKeyMUXOutput[5]), .B(
        AddKeyMUXOutput[7]), .Z(SubCellInst_LFInst_1_LFInst_2_n4 ) );
  AND2 SubCellInst_LFInst_1_LFInst_2_U5  ( .A(AddKeyMUXOutput[5]), .B(
        AddKeyMUXOutput[4]), .Z(SubCellInst_LFInst_1_LFInst_2_n6 ) );
  ORN2 SubCellInst_LFInst_1_LFInst_2_U4  ( .A(AddKeyMUXOutput[7]), .B(
        SubCellInst_LFInst_1_LFInst_2_n6 ), .Z(
        SubCellInst_LFInst_1_LFInst_2_n5 ) );
  AND2 SubCellInst_LFInst_1_LFInst_2_U3  ( .A(
        SubCellInst_LFInst_1_LFInst_2_n4 ), .B(
        SubCellInst_LFInst_1_LFInst_2_n5 ), .Z(
        SubCellInst_LFInst_1_LFInst_2_n3 ) );
  ORN2 SubCellInst_LFInst_1_LFInst_2_U2  ( .A(
        SubCellInst_LFInst_1_LFInst_2_n3 ), .B(AddKeyMUXOutput[6]), .Z(
        SubCellInst_LFInst_1_LFInst_2_n2 ) );
  ORN2 SubCellInst_LFInst_1_LFInst_2_U1  ( .A(
        SubCellInst_LFInst_1_LFInst_2_n1 ), .B(
        SubCellInst_LFInst_1_LFInst_2_n2 ), .Z(MCInst1_MC3_v3_0 [3]) );
  AND2 SubCellInst_LFInst_1_LFInst_1_U8  ( .A(AddKeyMUXOutput[6]), .B(
        AddKeyMUXOutput[4]), .Z(SubCellInst_LFInst_1_LFInst_1_n4 ) );
  AND2 SubCellInst_LFInst_1_LFInst_1_U7  ( .A(AddKeyMUXOutput[5]), .B(
        AddKeyMUXOutput[4]), .Z(SubCellInst_LFInst_1_LFInst_1_n7 ) );
  OR2 SubCellInst_LFInst_1_LFInst_1_U6  ( .A(AddKeyMUXOutput[6]), .B(
        SubCellInst_LFInst_1_LFInst_1_n7 ), .Z(
        SubCellInst_LFInst_1_LFInst_1_n6 ) );
  ORN2 SubCellInst_LFInst_1_LFInst_1_U5  ( .A(
        SubCellInst_LFInst_1_LFInst_1_n4 ), .B(
        SubCellInst_LFInst_1_LFInst_1_n6 ), .Z(
        SubCellInst_LFInst_1_LFInst_1_n5 ) );
  AND2 SubCellInst_LFInst_1_LFInst_1_U4  ( .A(AddKeyMUXOutput[7]), .B(
        SubCellInst_LFInst_1_LFInst_1_n5 ), .Z(
        SubCellInst_LFInst_1_LFInst_1_n1 ) );
  BIC2 SubCellInst_LFInst_1_LFInst_1_U3  ( .A(AddKeyMUXOutput[5]), .B(
        SubCellInst_LFInst_1_LFInst_1_n4 ), .Z(
        SubCellInst_LFInst_1_LFInst_1_n3 ) );
  ORN2 SubCellInst_LFInst_1_LFInst_1_U2  ( .A(AddKeyMUXOutput[7]), .B(
        SubCellInst_LFInst_1_LFInst_1_n3 ), .Z(
        SubCellInst_LFInst_1_LFInst_1_n2 ) );
  ORN2 SubCellInst_LFInst_1_LFInst_1_U1  ( .A(
        SubCellInst_LFInst_1_LFInst_1_n1 ), .B(
        SubCellInst_LFInst_1_LFInst_1_n2 ), .Z(MCInst1_MC3_v3_0 [2]) );
  BIC2 SubCellInst_LFInst_1_LFInst_0_U3  ( .A(AddKeyMUXOutput[6]), .B(
        AddKeyMUXOutput[5]), .Z(SubCellInst_LFInst_1_LFInst_0_n1 ) );
  XOR2 SubCellInst_LFInst_1_LFInst_0_U2  ( .A(AddKeyMUXOutput[7]), .B(
        AddKeyMUXOutput[4]), .Z(SubCellInst_LFInst_1_LFInst_0_n2 ) );
  XOR2 SubCellInst_LFInst_1_LFInst_0_U1  ( .A(
        SubCellInst_LFInst_1_LFInst_0_n1 ), .B(
        SubCellInst_LFInst_1_LFInst_0_n2 ), .Z(MCInst1_MC3_v3_2 [3]) );
  OR2 SubCellInst_LFInst_2_LFInst_3_U9  ( .A(AddConstOutput[1]), .B(
        AddConstOutput[0]), .Z(SubCellInst_LFInst_2_LFInst_3_n5 ) );
  AND2 SubCellInst_LFInst_2_LFInst_3_U8  ( .A(AddConstOutput[3]), .B(
        SubCellInst_LFInst_2_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_2_LFInst_3_n7 ) );
  AND2 SubCellInst_LFInst_2_LFInst_3_U7  ( .A(AddConstOutput[0]), .B(
        AddConstOutput[1]), .Z(SubCellInst_LFInst_2_LFInst_3_n8 ) );
  OR2 SubCellInst_LFInst_2_LFInst_3_U6  ( .A(
        SubCellInst_LFInst_2_LFInst_3_n7 ), .B(
        SubCellInst_LFInst_2_LFInst_3_n8 ), .Z(
        SubCellInst_LFInst_2_LFInst_3_n6 ) );
  BIC2 SubCellInst_LFInst_2_LFInst_3_U5  ( .A(
        SubCellInst_LFInst_2_LFInst_3_n6 ), .B(AddConstOutput[2]), .Z(
        SubCellInst_LFInst_2_LFInst_3_n1 ) );
  AND2 SubCellInst_LFInst_2_LFInst_3_U4  ( .A(AddConstOutput[2]), .B(
        AddConstOutput[1]), .Z(SubCellInst_LFInst_2_LFInst_3_n4 ) );
  ORN2 SubCellInst_LFInst_2_LFInst_3_U3  ( .A(
        SubCellInst_LFInst_2_LFInst_3_n4 ), .B(
        SubCellInst_LFInst_2_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_2_LFInst_3_n3 ) );
  ORN2 SubCellInst_LFInst_2_LFInst_3_U2  ( .A(AddConstOutput[3]), .B(
        SubCellInst_LFInst_2_LFInst_3_n3 ), .Z(
        SubCellInst_LFInst_2_LFInst_3_n2 ) );
  ORN2 SubCellInst_LFInst_2_LFInst_3_U1  ( .A(
        SubCellInst_LFInst_2_LFInst_3_n1 ), .B(
        SubCellInst_LFInst_2_LFInst_3_n2 ), .Z(MCInst1_MC2_v3_2 [2]) );
  BIC2 SubCellInst_LFInst_2_LFInst_2_U11  ( .A(AddConstOutput[1]), .B(
        AddConstOutput[0]), .Z(SubCellInst_LFInst_2_LFInst_2_n8 ) );
  ORN2 SubCellInst_LFInst_2_LFInst_2_U10  ( .A(AddConstOutput[0]), .B(
        AddConstOutput[3]), .Z(SubCellInst_LFInst_2_LFInst_2_n10 ) );
  ORN2 SubCellInst_LFInst_2_LFInst_2_U9  ( .A(AddConstOutput[1]), .B(
        SubCellInst_LFInst_2_LFInst_2_n10 ), .Z(
        SubCellInst_LFInst_2_LFInst_2_n9 ) );
  ORN2 SubCellInst_LFInst_2_LFInst_2_U8  ( .A(
        SubCellInst_LFInst_2_LFInst_2_n8 ), .B(
        SubCellInst_LFInst_2_LFInst_2_n9 ), .Z(
        SubCellInst_LFInst_2_LFInst_2_n7 ) );
  BIC2 SubCellInst_LFInst_2_LFInst_2_U7  ( .A(
        SubCellInst_LFInst_2_LFInst_2_n7 ), .B(AddConstOutput[2]), .Z(
        SubCellInst_LFInst_2_LFInst_2_n1 ) );
  ORN2 SubCellInst_LFInst_2_LFInst_2_U6  ( .A(AddConstOutput[1]), .B(
        AddConstOutput[3]), .Z(SubCellInst_LFInst_2_LFInst_2_n4 ) );
  AND2 SubCellInst_LFInst_2_LFInst_2_U5  ( .A(AddConstOutput[1]), .B(
        AddConstOutput[0]), .Z(SubCellInst_LFInst_2_LFInst_2_n6 ) );
  ORN2 SubCellInst_LFInst_2_LFInst_2_U4  ( .A(AddConstOutput[3]), .B(
        SubCellInst_LFInst_2_LFInst_2_n6 ), .Z(
        SubCellInst_LFInst_2_LFInst_2_n5 ) );
  AND2 SubCellInst_LFInst_2_LFInst_2_U3  ( .A(
        SubCellInst_LFInst_2_LFInst_2_n4 ), .B(
        SubCellInst_LFInst_2_LFInst_2_n5 ), .Z(
        SubCellInst_LFInst_2_LFInst_2_n3 ) );
  ORN2 SubCellInst_LFInst_2_LFInst_2_U2  ( .A(
        SubCellInst_LFInst_2_LFInst_2_n3 ), .B(AddConstOutput[2]), .Z(
        SubCellInst_LFInst_2_LFInst_2_n2 ) );
  ORN2 SubCellInst_LFInst_2_LFInst_2_U1  ( .A(
        SubCellInst_LFInst_2_LFInst_2_n1 ), .B(
        SubCellInst_LFInst_2_LFInst_2_n2 ), .Z(MCInst1_MC2_v3_0 [3]) );
  AND2 SubCellInst_LFInst_2_LFInst_1_U8  ( .A(AddConstOutput[2]), .B(
        AddConstOutput[0]), .Z(SubCellInst_LFInst_2_LFInst_1_n4 ) );
  AND2 SubCellInst_LFInst_2_LFInst_1_U7  ( .A(AddConstOutput[1]), .B(
        AddConstOutput[0]), .Z(SubCellInst_LFInst_2_LFInst_1_n7 ) );
  OR2 SubCellInst_LFInst_2_LFInst_1_U6  ( .A(AddConstOutput[2]), .B(
        SubCellInst_LFInst_2_LFInst_1_n7 ), .Z(
        SubCellInst_LFInst_2_LFInst_1_n6 ) );
  ORN2 SubCellInst_LFInst_2_LFInst_1_U5  ( .A(
        SubCellInst_LFInst_2_LFInst_1_n4 ), .B(
        SubCellInst_LFInst_2_LFInst_1_n6 ), .Z(
        SubCellInst_LFInst_2_LFInst_1_n5 ) );
  AND2 SubCellInst_LFInst_2_LFInst_1_U4  ( .A(AddConstOutput[3]), .B(
        SubCellInst_LFInst_2_LFInst_1_n5 ), .Z(
        SubCellInst_LFInst_2_LFInst_1_n1 ) );
  BIC2 SubCellInst_LFInst_2_LFInst_1_U3  ( .A(AddConstOutput[1]), .B(
        SubCellInst_LFInst_2_LFInst_1_n4 ), .Z(
        SubCellInst_LFInst_2_LFInst_1_n3 ) );
  ORN2 SubCellInst_LFInst_2_LFInst_1_U2  ( .A(AddConstOutput[3]), .B(
        SubCellInst_LFInst_2_LFInst_1_n3 ), .Z(
        SubCellInst_LFInst_2_LFInst_1_n2 ) );
  ORN2 SubCellInst_LFInst_2_LFInst_1_U1  ( .A(
        SubCellInst_LFInst_2_LFInst_1_n1 ), .B(
        SubCellInst_LFInst_2_LFInst_1_n2 ), .Z(MCInst1_MC2_v3_0 [2]) );
  BIC2 SubCellInst_LFInst_2_LFInst_0_U3  ( .A(AddConstOutput[2]), .B(
        AddConstOutput[1]), .Z(SubCellInst_LFInst_2_LFInst_0_n1 ) );
  XOR2 SubCellInst_LFInst_2_LFInst_0_U2  ( .A(AddConstOutput[3]), .B(
        AddConstOutput[0]), .Z(SubCellInst_LFInst_2_LFInst_0_n2 ) );
  XOR2 SubCellInst_LFInst_2_LFInst_0_U1  ( .A(
        SubCellInst_LFInst_2_LFInst_0_n1 ), .B(
        SubCellInst_LFInst_2_LFInst_0_n2 ), .Z(MCInst1_MC2_v3_2 [3]) );
  OR2 SubCellInst_LFInst_3_LFInst_3_U9  ( .A(AddConstOutput[5]), .B(
        AddConstOutput[4]), .Z(SubCellInst_LFInst_3_LFInst_3_n5 ) );
  AND2 SubCellInst_LFInst_3_LFInst_3_U8  ( .A(AddConstOutput[7]), .B(
        SubCellInst_LFInst_3_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_3_LFInst_3_n7 ) );
  AND2 SubCellInst_LFInst_3_LFInst_3_U7  ( .A(AddConstOutput[4]), .B(
        AddConstOutput[5]), .Z(SubCellInst_LFInst_3_LFInst_3_n8 ) );
  OR2 SubCellInst_LFInst_3_LFInst_3_U6  ( .A(
        SubCellInst_LFInst_3_LFInst_3_n7 ), .B(
        SubCellInst_LFInst_3_LFInst_3_n8 ), .Z(
        SubCellInst_LFInst_3_LFInst_3_n6 ) );
  BIC2 SubCellInst_LFInst_3_LFInst_3_U5  ( .A(
        SubCellInst_LFInst_3_LFInst_3_n6 ), .B(AddConstOutput[6]), .Z(
        SubCellInst_LFInst_3_LFInst_3_n1 ) );
  AND2 SubCellInst_LFInst_3_LFInst_3_U4  ( .A(AddConstOutput[6]), .B(
        AddConstOutput[5]), .Z(SubCellInst_LFInst_3_LFInst_3_n4 ) );
  ORN2 SubCellInst_LFInst_3_LFInst_3_U3  ( .A(
        SubCellInst_LFInst_3_LFInst_3_n4 ), .B(
        SubCellInst_LFInst_3_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_3_LFInst_3_n3 ) );
  ORN2 SubCellInst_LFInst_3_LFInst_3_U2  ( .A(AddConstOutput[7]), .B(
        SubCellInst_LFInst_3_LFInst_3_n3 ), .Z(
        SubCellInst_LFInst_3_LFInst_3_n2 ) );
  ORN2 SubCellInst_LFInst_3_LFInst_3_U1  ( .A(
        SubCellInst_LFInst_3_LFInst_3_n1 ), .B(
        SubCellInst_LFInst_3_LFInst_3_n2 ), .Z(MCInst1_MC1_v3_2 [2]) );
  BIC2 SubCellInst_LFInst_3_LFInst_2_U11  ( .A(AddConstOutput[5]), .B(
        AddConstOutput[4]), .Z(SubCellInst_LFInst_3_LFInst_2_n8 ) );
  ORN2 SubCellInst_LFInst_3_LFInst_2_U10  ( .A(AddConstOutput[4]), .B(
        AddConstOutput[7]), .Z(SubCellInst_LFInst_3_LFInst_2_n10 ) );
  ORN2 SubCellInst_LFInst_3_LFInst_2_U9  ( .A(AddConstOutput[5]), .B(
        SubCellInst_LFInst_3_LFInst_2_n10 ), .Z(
        SubCellInst_LFInst_3_LFInst_2_n9 ) );
  ORN2 SubCellInst_LFInst_3_LFInst_2_U8  ( .A(
        SubCellInst_LFInst_3_LFInst_2_n8 ), .B(
        SubCellInst_LFInst_3_LFInst_2_n9 ), .Z(
        SubCellInst_LFInst_3_LFInst_2_n7 ) );
  BIC2 SubCellInst_LFInst_3_LFInst_2_U7  ( .A(
        SubCellInst_LFInst_3_LFInst_2_n7 ), .B(AddConstOutput[6]), .Z(
        SubCellInst_LFInst_3_LFInst_2_n1 ) );
  ORN2 SubCellInst_LFInst_3_LFInst_2_U6  ( .A(AddConstOutput[5]), .B(
        AddConstOutput[7]), .Z(SubCellInst_LFInst_3_LFInst_2_n4 ) );
  AND2 SubCellInst_LFInst_3_LFInst_2_U5  ( .A(AddConstOutput[5]), .B(
        AddConstOutput[4]), .Z(SubCellInst_LFInst_3_LFInst_2_n6 ) );
  ORN2 SubCellInst_LFInst_3_LFInst_2_U4  ( .A(AddConstOutput[7]), .B(
        SubCellInst_LFInst_3_LFInst_2_n6 ), .Z(
        SubCellInst_LFInst_3_LFInst_2_n5 ) );
  AND2 SubCellInst_LFInst_3_LFInst_2_U3  ( .A(
        SubCellInst_LFInst_3_LFInst_2_n4 ), .B(
        SubCellInst_LFInst_3_LFInst_2_n5 ), .Z(
        SubCellInst_LFInst_3_LFInst_2_n3 ) );
  ORN2 SubCellInst_LFInst_3_LFInst_2_U2  ( .A(
        SubCellInst_LFInst_3_LFInst_2_n3 ), .B(AddConstOutput[6]), .Z(
        SubCellInst_LFInst_3_LFInst_2_n2 ) );
  ORN2 SubCellInst_LFInst_3_LFInst_2_U1  ( .A(
        SubCellInst_LFInst_3_LFInst_2_n1 ), .B(
        SubCellInst_LFInst_3_LFInst_2_n2 ), .Z(MCInst1_MC1_v3_0 [3]) );
  AND2 SubCellInst_LFInst_3_LFInst_1_U8  ( .A(AddConstOutput[6]), .B(
        AddConstOutput[4]), .Z(SubCellInst_LFInst_3_LFInst_1_n4 ) );
  AND2 SubCellInst_LFInst_3_LFInst_1_U7  ( .A(AddConstOutput[5]), .B(
        AddConstOutput[4]), .Z(SubCellInst_LFInst_3_LFInst_1_n7 ) );
  OR2 SubCellInst_LFInst_3_LFInst_1_U6  ( .A(AddConstOutput[6]), .B(
        SubCellInst_LFInst_3_LFInst_1_n7 ), .Z(
        SubCellInst_LFInst_3_LFInst_1_n6 ) );
  ORN2 SubCellInst_LFInst_3_LFInst_1_U5  ( .A(
        SubCellInst_LFInst_3_LFInst_1_n4 ), .B(
        SubCellInst_LFInst_3_LFInst_1_n6 ), .Z(
        SubCellInst_LFInst_3_LFInst_1_n5 ) );
  AND2 SubCellInst_LFInst_3_LFInst_1_U4  ( .A(AddConstOutput[7]), .B(
        SubCellInst_LFInst_3_LFInst_1_n5 ), .Z(
        SubCellInst_LFInst_3_LFInst_1_n1 ) );
  BIC2 SubCellInst_LFInst_3_LFInst_1_U3  ( .A(AddConstOutput[5]), .B(
        SubCellInst_LFInst_3_LFInst_1_n4 ), .Z(
        SubCellInst_LFInst_3_LFInst_1_n3 ) );
  ORN2 SubCellInst_LFInst_3_LFInst_1_U2  ( .A(AddConstOutput[7]), .B(
        SubCellInst_LFInst_3_LFInst_1_n3 ), .Z(
        SubCellInst_LFInst_3_LFInst_1_n2 ) );
  ORN2 SubCellInst_LFInst_3_LFInst_1_U1  ( .A(
        SubCellInst_LFInst_3_LFInst_1_n1 ), .B(
        SubCellInst_LFInst_3_LFInst_1_n2 ), .Z(MCInst1_MC1_v3_0 [2]) );
  BIC2 SubCellInst_LFInst_3_LFInst_0_U3  ( .A(AddConstOutput[6]), .B(
        AddConstOutput[5]), .Z(SubCellInst_LFInst_3_LFInst_0_n1 ) );
  XOR2 SubCellInst_LFInst_3_LFInst_0_U2  ( .A(AddConstOutput[7]), .B(
        AddConstOutput[4]), .Z(SubCellInst_LFInst_3_LFInst_0_n2 ) );
  XOR2 SubCellInst_LFInst_3_LFInst_0_U1  ( .A(
        SubCellInst_LFInst_3_LFInst_0_n1 ), .B(
        SubCellInst_LFInst_3_LFInst_0_n2 ), .Z(MCInst1_MC1_v3_2 [3]) );
  OR2 SubCellInst_LFInst_4_LFInst_3_U9  ( .A(AddKeyMUXOutput[17]), .B(
        AddKeyMUXOutput[16]), .Z(SubCellInst_LFInst_4_LFInst_3_n5 ) );
  AND2 SubCellInst_LFInst_4_LFInst_3_U8  ( .A(AddKeyMUXOutput[19]), .B(
        SubCellInst_LFInst_4_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_4_LFInst_3_n7 ) );
  AND2 SubCellInst_LFInst_4_LFInst_3_U7  ( .A(AddKeyMUXOutput[16]), .B(
        AddKeyMUXOutput[17]), .Z(SubCellInst_LFInst_4_LFInst_3_n8 ) );
  OR2 SubCellInst_LFInst_4_LFInst_3_U6  ( .A(
        SubCellInst_LFInst_4_LFInst_3_n7 ), .B(
        SubCellInst_LFInst_4_LFInst_3_n8 ), .Z(
        SubCellInst_LFInst_4_LFInst_3_n6 ) );
  BIC2 SubCellInst_LFInst_4_LFInst_3_U5  ( .A(
        SubCellInst_LFInst_4_LFInst_3_n6 ), .B(AddKeyMUXOutput[18]), .Z(
        SubCellInst_LFInst_4_LFInst_3_n1 ) );
  AND2 SubCellInst_LFInst_4_LFInst_3_U4  ( .A(AddKeyMUXOutput[18]), .B(
        AddKeyMUXOutput[17]), .Z(SubCellInst_LFInst_4_LFInst_3_n4 ) );
  ORN2 SubCellInst_LFInst_4_LFInst_3_U3  ( .A(
        SubCellInst_LFInst_4_LFInst_3_n4 ), .B(
        SubCellInst_LFInst_4_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_4_LFInst_3_n3 ) );
  ORN2 SubCellInst_LFInst_4_LFInst_3_U2  ( .A(AddKeyMUXOutput[19]), .B(
        SubCellInst_LFInst_4_LFInst_3_n3 ), .Z(
        SubCellInst_LFInst_4_LFInst_3_n2 ) );
  ORN2 SubCellInst_LFInst_4_LFInst_3_U1  ( .A(
        SubCellInst_LFInst_4_LFInst_3_n1 ), .B(
        SubCellInst_LFInst_4_LFInst_3_n2 ), .Z(MCInst1_MC1_v2_0 [0]) );
  BIC2 SubCellInst_LFInst_4_LFInst_2_U11  ( .A(AddKeyMUXOutput[17]), .B(
        AddKeyMUXOutput[16]), .Z(SubCellInst_LFInst_4_LFInst_2_n8 ) );
  ORN2 SubCellInst_LFInst_4_LFInst_2_U10  ( .A(AddKeyMUXOutput[16]), .B(
        AddKeyMUXOutput[19]), .Z(SubCellInst_LFInst_4_LFInst_2_n10 ) );
  ORN2 SubCellInst_LFInst_4_LFInst_2_U9  ( .A(AddKeyMUXOutput[17]), .B(
        SubCellInst_LFInst_4_LFInst_2_n10 ), .Z(
        SubCellInst_LFInst_4_LFInst_2_n9 ) );
  ORN2 SubCellInst_LFInst_4_LFInst_2_U8  ( .A(
        SubCellInst_LFInst_4_LFInst_2_n8 ), .B(
        SubCellInst_LFInst_4_LFInst_2_n9 ), .Z(
        SubCellInst_LFInst_4_LFInst_2_n7 ) );
  BIC2 SubCellInst_LFInst_4_LFInst_2_U7  ( .A(
        SubCellInst_LFInst_4_LFInst_2_n7 ), .B(AddKeyMUXOutput[18]), .Z(
        SubCellInst_LFInst_4_LFInst_2_n1 ) );
  ORN2 SubCellInst_LFInst_4_LFInst_2_U6  ( .A(AddKeyMUXOutput[17]), .B(
        AddKeyMUXOutput[19]), .Z(SubCellInst_LFInst_4_LFInst_2_n4 ) );
  AND2 SubCellInst_LFInst_4_LFInst_2_U5  ( .A(AddKeyMUXOutput[17]), .B(
        AddKeyMUXOutput[16]), .Z(SubCellInst_LFInst_4_LFInst_2_n6 ) );
  ORN2 SubCellInst_LFInst_4_LFInst_2_U4  ( .A(AddKeyMUXOutput[19]), .B(
        SubCellInst_LFInst_4_LFInst_2_n6 ), .Z(
        SubCellInst_LFInst_4_LFInst_2_n5 ) );
  AND2 SubCellInst_LFInst_4_LFInst_2_U3  ( .A(
        SubCellInst_LFInst_4_LFInst_2_n4 ), .B(
        SubCellInst_LFInst_4_LFInst_2_n5 ), .Z(
        SubCellInst_LFInst_4_LFInst_2_n3 ) );
  ORN2 SubCellInst_LFInst_4_LFInst_2_U2  ( .A(
        SubCellInst_LFInst_4_LFInst_2_n3 ), .B(AddKeyMUXOutput[18]), .Z(
        SubCellInst_LFInst_4_LFInst_2_n2 ) );
  ORN2 SubCellInst_LFInst_4_LFInst_2_U1  ( .A(
        SubCellInst_LFInst_4_LFInst_2_n1 ), .B(
        SubCellInst_LFInst_4_LFInst_2_n2 ), .Z(MCInst1_MC1_v2_0 [3]) );
  AND2 SubCellInst_LFInst_4_LFInst_1_U8  ( .A(AddKeyMUXOutput[18]), .B(
        AddKeyMUXOutput[16]), .Z(SubCellInst_LFInst_4_LFInst_1_n4 ) );
  AND2 SubCellInst_LFInst_4_LFInst_1_U7  ( .A(AddKeyMUXOutput[17]), .B(
        AddKeyMUXOutput[16]), .Z(SubCellInst_LFInst_4_LFInst_1_n7 ) );
  OR2 SubCellInst_LFInst_4_LFInst_1_U6  ( .A(AddKeyMUXOutput[18]), .B(
        SubCellInst_LFInst_4_LFInst_1_n7 ), .Z(
        SubCellInst_LFInst_4_LFInst_1_n6 ) );
  ORN2 SubCellInst_LFInst_4_LFInst_1_U5  ( .A(
        SubCellInst_LFInst_4_LFInst_1_n4 ), .B(
        SubCellInst_LFInst_4_LFInst_1_n6 ), .Z(
        SubCellInst_LFInst_4_LFInst_1_n5 ) );
  AND2 SubCellInst_LFInst_4_LFInst_1_U4  ( .A(AddKeyMUXOutput[19]), .B(
        SubCellInst_LFInst_4_LFInst_1_n5 ), .Z(
        SubCellInst_LFInst_4_LFInst_1_n1 ) );
  BIC2 SubCellInst_LFInst_4_LFInst_1_U3  ( .A(AddKeyMUXOutput[17]), .B(
        SubCellInst_LFInst_4_LFInst_1_n4 ), .Z(
        SubCellInst_LFInst_4_LFInst_1_n3 ) );
  ORN2 SubCellInst_LFInst_4_LFInst_1_U2  ( .A(AddKeyMUXOutput[19]), .B(
        SubCellInst_LFInst_4_LFInst_1_n3 ), .Z(
        SubCellInst_LFInst_4_LFInst_1_n2 ) );
  ORN2 SubCellInst_LFInst_4_LFInst_1_U1  ( .A(
        SubCellInst_LFInst_4_LFInst_1_n1 ), .B(
        SubCellInst_LFInst_4_LFInst_1_n2 ), .Z(MCInst1_MC1_v2_0 [2]) );
  BIC2 SubCellInst_LFInst_4_LFInst_0_U3  ( .A(AddKeyMUXOutput[18]), .B(
        AddKeyMUXOutput[17]), .Z(SubCellInst_LFInst_4_LFInst_0_n1 ) );
  XOR2 SubCellInst_LFInst_4_LFInst_0_U2  ( .A(AddKeyMUXOutput[19]), .B(
        AddKeyMUXOutput[16]), .Z(SubCellInst_LFInst_4_LFInst_0_n2 ) );
  XOR2 SubCellInst_LFInst_4_LFInst_0_U1  ( .A(
        SubCellInst_LFInst_4_LFInst_0_n1 ), .B(
        SubCellInst_LFInst_4_LFInst_0_n2 ), .Z(MCInst1_MC1_v2_3 [1]) );
  OR2 SubCellInst_LFInst_5_LFInst_3_U9  ( .A(AddKeyMUXOutput[21]), .B(
        AddKeyMUXOutput[20]), .Z(SubCellInst_LFInst_5_LFInst_3_n5 ) );
  AND2 SubCellInst_LFInst_5_LFInst_3_U8  ( .A(AddKeyMUXOutput[23]), .B(
        SubCellInst_LFInst_5_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_5_LFInst_3_n7 ) );
  AND2 SubCellInst_LFInst_5_LFInst_3_U7  ( .A(AddKeyMUXOutput[20]), .B(
        AddKeyMUXOutput[21]), .Z(SubCellInst_LFInst_5_LFInst_3_n8 ) );
  OR2 SubCellInst_LFInst_5_LFInst_3_U6  ( .A(
        SubCellInst_LFInst_5_LFInst_3_n7 ), .B(
        SubCellInst_LFInst_5_LFInst_3_n8 ), .Z(
        SubCellInst_LFInst_5_LFInst_3_n6 ) );
  BIC2 SubCellInst_LFInst_5_LFInst_3_U5  ( .A(
        SubCellInst_LFInst_5_LFInst_3_n6 ), .B(AddKeyMUXOutput[22]), .Z(
        SubCellInst_LFInst_5_LFInst_3_n1 ) );
  AND2 SubCellInst_LFInst_5_LFInst_3_U4  ( .A(AddKeyMUXOutput[22]), .B(
        AddKeyMUXOutput[21]), .Z(SubCellInst_LFInst_5_LFInst_3_n4 ) );
  ORN2 SubCellInst_LFInst_5_LFInst_3_U3  ( .A(
        SubCellInst_LFInst_5_LFInst_3_n4 ), .B(
        SubCellInst_LFInst_5_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_5_LFInst_3_n3 ) );
  ORN2 SubCellInst_LFInst_5_LFInst_3_U2  ( .A(AddKeyMUXOutput[23]), .B(
        SubCellInst_LFInst_5_LFInst_3_n3 ), .Z(
        SubCellInst_LFInst_5_LFInst_3_n2 ) );
  ORN2 SubCellInst_LFInst_5_LFInst_3_U1  ( .A(
        SubCellInst_LFInst_5_LFInst_3_n1 ), .B(
        SubCellInst_LFInst_5_LFInst_3_n2 ), .Z(MCInst1_MC0_v2_0 [0]) );
  BIC2 SubCellInst_LFInst_5_LFInst_2_U11  ( .A(AddKeyMUXOutput[21]), .B(
        AddKeyMUXOutput[20]), .Z(SubCellInst_LFInst_5_LFInst_2_n8 ) );
  ORN2 SubCellInst_LFInst_5_LFInst_2_U10  ( .A(AddKeyMUXOutput[20]), .B(
        AddKeyMUXOutput[23]), .Z(SubCellInst_LFInst_5_LFInst_2_n10 ) );
  ORN2 SubCellInst_LFInst_5_LFInst_2_U9  ( .A(AddKeyMUXOutput[21]), .B(
        SubCellInst_LFInst_5_LFInst_2_n10 ), .Z(
        SubCellInst_LFInst_5_LFInst_2_n9 ) );
  ORN2 SubCellInst_LFInst_5_LFInst_2_U8  ( .A(
        SubCellInst_LFInst_5_LFInst_2_n8 ), .B(
        SubCellInst_LFInst_5_LFInst_2_n9 ), .Z(
        SubCellInst_LFInst_5_LFInst_2_n7 ) );
  BIC2 SubCellInst_LFInst_5_LFInst_2_U7  ( .A(
        SubCellInst_LFInst_5_LFInst_2_n7 ), .B(AddKeyMUXOutput[22]), .Z(
        SubCellInst_LFInst_5_LFInst_2_n1 ) );
  ORN2 SubCellInst_LFInst_5_LFInst_2_U6  ( .A(AddKeyMUXOutput[21]), .B(
        AddKeyMUXOutput[23]), .Z(SubCellInst_LFInst_5_LFInst_2_n4 ) );
  AND2 SubCellInst_LFInst_5_LFInst_2_U5  ( .A(AddKeyMUXOutput[21]), .B(
        AddKeyMUXOutput[20]), .Z(SubCellInst_LFInst_5_LFInst_2_n6 ) );
  ORN2 SubCellInst_LFInst_5_LFInst_2_U4  ( .A(AddKeyMUXOutput[23]), .B(
        SubCellInst_LFInst_5_LFInst_2_n6 ), .Z(
        SubCellInst_LFInst_5_LFInst_2_n5 ) );
  AND2 SubCellInst_LFInst_5_LFInst_2_U3  ( .A(
        SubCellInst_LFInst_5_LFInst_2_n4 ), .B(
        SubCellInst_LFInst_5_LFInst_2_n5 ), .Z(
        SubCellInst_LFInst_5_LFInst_2_n3 ) );
  ORN2 SubCellInst_LFInst_5_LFInst_2_U2  ( .A(
        SubCellInst_LFInst_5_LFInst_2_n3 ), .B(AddKeyMUXOutput[22]), .Z(
        SubCellInst_LFInst_5_LFInst_2_n2 ) );
  ORN2 SubCellInst_LFInst_5_LFInst_2_U1  ( .A(
        SubCellInst_LFInst_5_LFInst_2_n1 ), .B(
        SubCellInst_LFInst_5_LFInst_2_n2 ), .Z(MCInst1_MC0_v2_0 [3]) );
  AND2 SubCellInst_LFInst_5_LFInst_1_U8  ( .A(AddKeyMUXOutput[22]), .B(
        AddKeyMUXOutput[20]), .Z(SubCellInst_LFInst_5_LFInst_1_n4 ) );
  AND2 SubCellInst_LFInst_5_LFInst_1_U7  ( .A(AddKeyMUXOutput[21]), .B(
        AddKeyMUXOutput[20]), .Z(SubCellInst_LFInst_5_LFInst_1_n7 ) );
  OR2 SubCellInst_LFInst_5_LFInst_1_U6  ( .A(AddKeyMUXOutput[22]), .B(
        SubCellInst_LFInst_5_LFInst_1_n7 ), .Z(
        SubCellInst_LFInst_5_LFInst_1_n6 ) );
  ORN2 SubCellInst_LFInst_5_LFInst_1_U5  ( .A(
        SubCellInst_LFInst_5_LFInst_1_n4 ), .B(
        SubCellInst_LFInst_5_LFInst_1_n6 ), .Z(
        SubCellInst_LFInst_5_LFInst_1_n5 ) );
  AND2 SubCellInst_LFInst_5_LFInst_1_U4  ( .A(AddKeyMUXOutput[23]), .B(
        SubCellInst_LFInst_5_LFInst_1_n5 ), .Z(
        SubCellInst_LFInst_5_LFInst_1_n1 ) );
  BIC2 SubCellInst_LFInst_5_LFInst_1_U3  ( .A(AddKeyMUXOutput[21]), .B(
        SubCellInst_LFInst_5_LFInst_1_n4 ), .Z(
        SubCellInst_LFInst_5_LFInst_1_n3 ) );
  ORN2 SubCellInst_LFInst_5_LFInst_1_U2  ( .A(AddKeyMUXOutput[23]), .B(
        SubCellInst_LFInst_5_LFInst_1_n3 ), .Z(
        SubCellInst_LFInst_5_LFInst_1_n2 ) );
  ORN2 SubCellInst_LFInst_5_LFInst_1_U1  ( .A(
        SubCellInst_LFInst_5_LFInst_1_n1 ), .B(
        SubCellInst_LFInst_5_LFInst_1_n2 ), .Z(MCInst1_MC0_v2_0 [2]) );
  BIC2 SubCellInst_LFInst_5_LFInst_0_U3  ( .A(AddKeyMUXOutput[22]), .B(
        AddKeyMUXOutput[21]), .Z(SubCellInst_LFInst_5_LFInst_0_n1 ) );
  XOR2 SubCellInst_LFInst_5_LFInst_0_U2  ( .A(AddKeyMUXOutput[23]), .B(
        AddKeyMUXOutput[20]), .Z(SubCellInst_LFInst_5_LFInst_0_n2 ) );
  XOR2 SubCellInst_LFInst_5_LFInst_0_U1  ( .A(
        SubCellInst_LFInst_5_LFInst_0_n1 ), .B(
        SubCellInst_LFInst_5_LFInst_0_n2 ), .Z(MCInst1_MC0_v2_3 [1]) );
  OR2 SubCellInst_LFInst_6_LFInst_3_U9  ( .A(AddConstOutput[9]), .B(
        AddConstOutput[8]), .Z(SubCellInst_LFInst_6_LFInst_3_n5 ) );
  AND2 SubCellInst_LFInst_6_LFInst_3_U8  ( .A(AddConstOutput[11]), .B(
        SubCellInst_LFInst_6_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_6_LFInst_3_n7 ) );
  AND2 SubCellInst_LFInst_6_LFInst_3_U7  ( .A(AddConstOutput[8]), .B(
        AddConstOutput[9]), .Z(SubCellInst_LFInst_6_LFInst_3_n8 ) );
  OR2 SubCellInst_LFInst_6_LFInst_3_U6  ( .A(
        SubCellInst_LFInst_6_LFInst_3_n7 ), .B(
        SubCellInst_LFInst_6_LFInst_3_n8 ), .Z(
        SubCellInst_LFInst_6_LFInst_3_n6 ) );
  BIC2 SubCellInst_LFInst_6_LFInst_3_U5  ( .A(
        SubCellInst_LFInst_6_LFInst_3_n6 ), .B(AddConstOutput[10]), .Z(
        SubCellInst_LFInst_6_LFInst_3_n1 ) );
  AND2 SubCellInst_LFInst_6_LFInst_3_U4  ( .A(AddConstOutput[10]), .B(
        AddConstOutput[9]), .Z(SubCellInst_LFInst_6_LFInst_3_n4 ) );
  ORN2 SubCellInst_LFInst_6_LFInst_3_U3  ( .A(
        SubCellInst_LFInst_6_LFInst_3_n4 ), .B(
        SubCellInst_LFInst_6_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_6_LFInst_3_n3 ) );
  ORN2 SubCellInst_LFInst_6_LFInst_3_U2  ( .A(AddConstOutput[11]), .B(
        SubCellInst_LFInst_6_LFInst_3_n3 ), .Z(
        SubCellInst_LFInst_6_LFInst_3_n2 ) );
  ORN2 SubCellInst_LFInst_6_LFInst_3_U1  ( .A(
        SubCellInst_LFInst_6_LFInst_3_n1 ), .B(
        SubCellInst_LFInst_6_LFInst_3_n2 ), .Z(MCInst1_MC3_v2_0 [0]) );
  BIC2 SubCellInst_LFInst_6_LFInst_2_U11  ( .A(AddConstOutput[9]), .B(
        AddConstOutput[8]), .Z(SubCellInst_LFInst_6_LFInst_2_n8 ) );
  ORN2 SubCellInst_LFInst_6_LFInst_2_U10  ( .A(AddConstOutput[8]), .B(
        AddConstOutput[11]), .Z(SubCellInst_LFInst_6_LFInst_2_n10 ) );
  ORN2 SubCellInst_LFInst_6_LFInst_2_U9  ( .A(AddConstOutput[9]), .B(
        SubCellInst_LFInst_6_LFInst_2_n10 ), .Z(
        SubCellInst_LFInst_6_LFInst_2_n9 ) );
  ORN2 SubCellInst_LFInst_6_LFInst_2_U8  ( .A(
        SubCellInst_LFInst_6_LFInst_2_n8 ), .B(
        SubCellInst_LFInst_6_LFInst_2_n9 ), .Z(
        SubCellInst_LFInst_6_LFInst_2_n7 ) );
  BIC2 SubCellInst_LFInst_6_LFInst_2_U7  ( .A(
        SubCellInst_LFInst_6_LFInst_2_n7 ), .B(AddConstOutput[10]), .Z(
        SubCellInst_LFInst_6_LFInst_2_n1 ) );
  ORN2 SubCellInst_LFInst_6_LFInst_2_U6  ( .A(AddConstOutput[9]), .B(
        AddConstOutput[11]), .Z(SubCellInst_LFInst_6_LFInst_2_n4 ) );
  AND2 SubCellInst_LFInst_6_LFInst_2_U5  ( .A(AddConstOutput[9]), .B(
        AddConstOutput[8]), .Z(SubCellInst_LFInst_6_LFInst_2_n6 ) );
  ORN2 SubCellInst_LFInst_6_LFInst_2_U4  ( .A(AddConstOutput[11]), .B(
        SubCellInst_LFInst_6_LFInst_2_n6 ), .Z(
        SubCellInst_LFInst_6_LFInst_2_n5 ) );
  AND2 SubCellInst_LFInst_6_LFInst_2_U3  ( .A(
        SubCellInst_LFInst_6_LFInst_2_n4 ), .B(
        SubCellInst_LFInst_6_LFInst_2_n5 ), .Z(
        SubCellInst_LFInst_6_LFInst_2_n3 ) );
  ORN2 SubCellInst_LFInst_6_LFInst_2_U2  ( .A(
        SubCellInst_LFInst_6_LFInst_2_n3 ), .B(AddConstOutput[10]), .Z(
        SubCellInst_LFInst_6_LFInst_2_n2 ) );
  ORN2 SubCellInst_LFInst_6_LFInst_2_U1  ( .A(
        SubCellInst_LFInst_6_LFInst_2_n1 ), .B(
        SubCellInst_LFInst_6_LFInst_2_n2 ), .Z(MCInst1_MC3_v2_0 [3]) );
  AND2 SubCellInst_LFInst_6_LFInst_1_U8  ( .A(AddConstOutput[10]), .B(
        AddConstOutput[8]), .Z(SubCellInst_LFInst_6_LFInst_1_n4 ) );
  AND2 SubCellInst_LFInst_6_LFInst_1_U7  ( .A(AddConstOutput[9]), .B(
        AddConstOutput[8]), .Z(SubCellInst_LFInst_6_LFInst_1_n7 ) );
  OR2 SubCellInst_LFInst_6_LFInst_1_U6  ( .A(AddConstOutput[10]), .B(
        SubCellInst_LFInst_6_LFInst_1_n7 ), .Z(
        SubCellInst_LFInst_6_LFInst_1_n6 ) );
  ORN2 SubCellInst_LFInst_6_LFInst_1_U5  ( .A(
        SubCellInst_LFInst_6_LFInst_1_n4 ), .B(
        SubCellInst_LFInst_6_LFInst_1_n6 ), .Z(
        SubCellInst_LFInst_6_LFInst_1_n5 ) );
  AND2 SubCellInst_LFInst_6_LFInst_1_U4  ( .A(AddConstOutput[11]), .B(
        SubCellInst_LFInst_6_LFInst_1_n5 ), .Z(
        SubCellInst_LFInst_6_LFInst_1_n1 ) );
  BIC2 SubCellInst_LFInst_6_LFInst_1_U3  ( .A(AddConstOutput[9]), .B(
        SubCellInst_LFInst_6_LFInst_1_n4 ), .Z(
        SubCellInst_LFInst_6_LFInst_1_n3 ) );
  ORN2 SubCellInst_LFInst_6_LFInst_1_U2  ( .A(AddConstOutput[11]), .B(
        SubCellInst_LFInst_6_LFInst_1_n3 ), .Z(
        SubCellInst_LFInst_6_LFInst_1_n2 ) );
  ORN2 SubCellInst_LFInst_6_LFInst_1_U1  ( .A(
        SubCellInst_LFInst_6_LFInst_1_n1 ), .B(
        SubCellInst_LFInst_6_LFInst_1_n2 ), .Z(MCInst1_MC3_v2_0 [2]) );
  BIC2 SubCellInst_LFInst_6_LFInst_0_U3  ( .A(AddConstOutput[10]), .B(
        AddConstOutput[9]), .Z(SubCellInst_LFInst_6_LFInst_0_n1 ) );
  XOR2 SubCellInst_LFInst_6_LFInst_0_U2  ( .A(AddConstOutput[11]), .B(
        AddConstOutput[8]), .Z(SubCellInst_LFInst_6_LFInst_0_n2 ) );
  XOR2 SubCellInst_LFInst_6_LFInst_0_U1  ( .A(
        SubCellInst_LFInst_6_LFInst_0_n1 ), .B(
        SubCellInst_LFInst_6_LFInst_0_n2 ), .Z(MCInst1_MC3_v2_3 [1]) );
  OR2 SubCellInst_LFInst_7_LFInst_3_U9  ( .A(AddConstOutput[13]), .B(
        AddConstOutput[12]), .Z(SubCellInst_LFInst_7_LFInst_3_n5 ) );
  AND2 SubCellInst_LFInst_7_LFInst_3_U8  ( .A(AddConstOutput[15]), .B(
        SubCellInst_LFInst_7_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_7_LFInst_3_n7 ) );
  AND2 SubCellInst_LFInst_7_LFInst_3_U7  ( .A(AddConstOutput[12]), .B(
        AddConstOutput[13]), .Z(SubCellInst_LFInst_7_LFInst_3_n8 ) );
  OR2 SubCellInst_LFInst_7_LFInst_3_U6  ( .A(
        SubCellInst_LFInst_7_LFInst_3_n7 ), .B(
        SubCellInst_LFInst_7_LFInst_3_n8 ), .Z(
        SubCellInst_LFInst_7_LFInst_3_n6 ) );
  BIC2 SubCellInst_LFInst_7_LFInst_3_U5  ( .A(
        SubCellInst_LFInst_7_LFInst_3_n6 ), .B(AddConstOutput[14]), .Z(
        SubCellInst_LFInst_7_LFInst_3_n1 ) );
  AND2 SubCellInst_LFInst_7_LFInst_3_U4  ( .A(AddConstOutput[14]), .B(
        AddConstOutput[13]), .Z(SubCellInst_LFInst_7_LFInst_3_n4 ) );
  ORN2 SubCellInst_LFInst_7_LFInst_3_U3  ( .A(
        SubCellInst_LFInst_7_LFInst_3_n4 ), .B(
        SubCellInst_LFInst_7_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_7_LFInst_3_n3 ) );
  ORN2 SubCellInst_LFInst_7_LFInst_3_U2  ( .A(AddConstOutput[15]), .B(
        SubCellInst_LFInst_7_LFInst_3_n3 ), .Z(
        SubCellInst_LFInst_7_LFInst_3_n2 ) );
  ORN2 SubCellInst_LFInst_7_LFInst_3_U1  ( .A(
        SubCellInst_LFInst_7_LFInst_3_n1 ), .B(
        SubCellInst_LFInst_7_LFInst_3_n2 ), .Z(MCInst1_MC2_v2_0 [0]) );
  BIC2 SubCellInst_LFInst_7_LFInst_2_U11  ( .A(AddConstOutput[13]), .B(
        AddConstOutput[12]), .Z(SubCellInst_LFInst_7_LFInst_2_n8 ) );
  ORN2 SubCellInst_LFInst_7_LFInst_2_U10  ( .A(AddConstOutput[12]), .B(
        AddConstOutput[15]), .Z(SubCellInst_LFInst_7_LFInst_2_n10 ) );
  ORN2 SubCellInst_LFInst_7_LFInst_2_U9  ( .A(AddConstOutput[13]), .B(
        SubCellInst_LFInst_7_LFInst_2_n10 ), .Z(
        SubCellInst_LFInst_7_LFInst_2_n9 ) );
  ORN2 SubCellInst_LFInst_7_LFInst_2_U8  ( .A(
        SubCellInst_LFInst_7_LFInst_2_n8 ), .B(
        SubCellInst_LFInst_7_LFInst_2_n9 ), .Z(
        SubCellInst_LFInst_7_LFInst_2_n7 ) );
  BIC2 SubCellInst_LFInst_7_LFInst_2_U7  ( .A(
        SubCellInst_LFInst_7_LFInst_2_n7 ), .B(AddConstOutput[14]), .Z(
        SubCellInst_LFInst_7_LFInst_2_n1 ) );
  ORN2 SubCellInst_LFInst_7_LFInst_2_U6  ( .A(AddConstOutput[13]), .B(
        AddConstOutput[15]), .Z(SubCellInst_LFInst_7_LFInst_2_n4 ) );
  AND2 SubCellInst_LFInst_7_LFInst_2_U5  ( .A(AddConstOutput[13]), .B(
        AddConstOutput[12]), .Z(SubCellInst_LFInst_7_LFInst_2_n6 ) );
  ORN2 SubCellInst_LFInst_7_LFInst_2_U4  ( .A(AddConstOutput[15]), .B(
        SubCellInst_LFInst_7_LFInst_2_n6 ), .Z(
        SubCellInst_LFInst_7_LFInst_2_n5 ) );
  AND2 SubCellInst_LFInst_7_LFInst_2_U3  ( .A(
        SubCellInst_LFInst_7_LFInst_2_n4 ), .B(
        SubCellInst_LFInst_7_LFInst_2_n5 ), .Z(
        SubCellInst_LFInst_7_LFInst_2_n3 ) );
  ORN2 SubCellInst_LFInst_7_LFInst_2_U2  ( .A(
        SubCellInst_LFInst_7_LFInst_2_n3 ), .B(AddConstOutput[14]), .Z(
        SubCellInst_LFInst_7_LFInst_2_n2 ) );
  ORN2 SubCellInst_LFInst_7_LFInst_2_U1  ( .A(
        SubCellInst_LFInst_7_LFInst_2_n1 ), .B(
        SubCellInst_LFInst_7_LFInst_2_n2 ), .Z(MCInst1_MC2_v2_0 [3]) );
  AND2 SubCellInst_LFInst_7_LFInst_1_U8  ( .A(AddConstOutput[14]), .B(
        AddConstOutput[12]), .Z(SubCellInst_LFInst_7_LFInst_1_n4 ) );
  AND2 SubCellInst_LFInst_7_LFInst_1_U7  ( .A(AddConstOutput[13]), .B(
        AddConstOutput[12]), .Z(SubCellInst_LFInst_7_LFInst_1_n7 ) );
  OR2 SubCellInst_LFInst_7_LFInst_1_U6  ( .A(AddConstOutput[14]), .B(
        SubCellInst_LFInst_7_LFInst_1_n7 ), .Z(
        SubCellInst_LFInst_7_LFInst_1_n6 ) );
  ORN2 SubCellInst_LFInst_7_LFInst_1_U5  ( .A(
        SubCellInst_LFInst_7_LFInst_1_n4 ), .B(
        SubCellInst_LFInst_7_LFInst_1_n6 ), .Z(
        SubCellInst_LFInst_7_LFInst_1_n5 ) );
  AND2 SubCellInst_LFInst_7_LFInst_1_U4  ( .A(AddConstOutput[15]), .B(
        SubCellInst_LFInst_7_LFInst_1_n5 ), .Z(
        SubCellInst_LFInst_7_LFInst_1_n1 ) );
  BIC2 SubCellInst_LFInst_7_LFInst_1_U3  ( .A(AddConstOutput[13]), .B(
        SubCellInst_LFInst_7_LFInst_1_n4 ), .Z(
        SubCellInst_LFInst_7_LFInst_1_n3 ) );
  ORN2 SubCellInst_LFInst_7_LFInst_1_U2  ( .A(AddConstOutput[15]), .B(
        SubCellInst_LFInst_7_LFInst_1_n3 ), .Z(
        SubCellInst_LFInst_7_LFInst_1_n2 ) );
  ORN2 SubCellInst_LFInst_7_LFInst_1_U1  ( .A(
        SubCellInst_LFInst_7_LFInst_1_n1 ), .B(
        SubCellInst_LFInst_7_LFInst_1_n2 ), .Z(MCInst1_MC2_v2_0 [2]) );
  BIC2 SubCellInst_LFInst_7_LFInst_0_U3  ( .A(AddConstOutput[14]), .B(
        AddConstOutput[13]), .Z(SubCellInst_LFInst_7_LFInst_0_n1 ) );
  XOR2 SubCellInst_LFInst_7_LFInst_0_U2  ( .A(AddConstOutput[15]), .B(
        AddConstOutput[12]), .Z(SubCellInst_LFInst_7_LFInst_0_n2 ) );
  XOR2 SubCellInst_LFInst_7_LFInst_0_U1  ( .A(
        SubCellInst_LFInst_7_LFInst_0_n1 ), .B(
        SubCellInst_LFInst_7_LFInst_0_n2 ), .Z(MCInst1_MC2_v2_3 [1]) );
  OR2 SubCellInst_LFInst_8_LFInst_3_U9  ( .A(AddKeyMUXOutput[33]), .B(
        AddKeyMUXOutput[32]), .Z(SubCellInst_LFInst_8_LFInst_3_n5 ) );
  AND2 SubCellInst_LFInst_8_LFInst_3_U8  ( .A(AddKeyMUXOutput[35]), .B(
        SubCellInst_LFInst_8_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_8_LFInst_3_n7 ) );
  AND2 SubCellInst_LFInst_8_LFInst_3_U7  ( .A(AddKeyMUXOutput[32]), .B(
        AddKeyMUXOutput[33]), .Z(SubCellInst_LFInst_8_LFInst_3_n8 ) );
  OR2 SubCellInst_LFInst_8_LFInst_3_U6  ( .A(
        SubCellInst_LFInst_8_LFInst_3_n7 ), .B(
        SubCellInst_LFInst_8_LFInst_3_n8 ), .Z(
        SubCellInst_LFInst_8_LFInst_3_n6 ) );
  BIC2 SubCellInst_LFInst_8_LFInst_3_U5  ( .A(
        SubCellInst_LFInst_8_LFInst_3_n6 ), .B(AddKeyMUXOutput[34]), .Z(
        SubCellInst_LFInst_8_LFInst_3_n1 ) );
  AND2 SubCellInst_LFInst_8_LFInst_3_U4  ( .A(AddKeyMUXOutput[34]), .B(
        AddKeyMUXOutput[33]), .Z(SubCellInst_LFInst_8_LFInst_3_n4 ) );
  ORN2 SubCellInst_LFInst_8_LFInst_3_U3  ( .A(
        SubCellInst_LFInst_8_LFInst_3_n4 ), .B(
        SubCellInst_LFInst_8_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_8_LFInst_3_n3 ) );
  ORN2 SubCellInst_LFInst_8_LFInst_3_U2  ( .A(AddKeyMUXOutput[35]), .B(
        SubCellInst_LFInst_8_LFInst_3_n3 ), .Z(
        SubCellInst_LFInst_8_LFInst_3_n2 ) );
  ORN2 SubCellInst_LFInst_8_LFInst_3_U1  ( .A(
        SubCellInst_LFInst_8_LFInst_3_n1 ), .B(
        SubCellInst_LFInst_8_LFInst_3_n2 ), .Z(MCInst1_MC2_v1_3 [0]) );
  BIC2 SubCellInst_LFInst_8_LFInst_2_U11  ( .A(AddKeyMUXOutput[33]), .B(
        AddKeyMUXOutput[32]), .Z(SubCellInst_LFInst_8_LFInst_2_n8 ) );
  ORN2 SubCellInst_LFInst_8_LFInst_2_U10  ( .A(AddKeyMUXOutput[32]), .B(
        AddKeyMUXOutput[35]), .Z(SubCellInst_LFInst_8_LFInst_2_n10 ) );
  ORN2 SubCellInst_LFInst_8_LFInst_2_U9  ( .A(AddKeyMUXOutput[33]), .B(
        SubCellInst_LFInst_8_LFInst_2_n10 ), .Z(
        SubCellInst_LFInst_8_LFInst_2_n9 ) );
  ORN2 SubCellInst_LFInst_8_LFInst_2_U8  ( .A(
        SubCellInst_LFInst_8_LFInst_2_n8 ), .B(
        SubCellInst_LFInst_8_LFInst_2_n9 ), .Z(
        SubCellInst_LFInst_8_LFInst_2_n7 ) );
  BIC2 SubCellInst_LFInst_8_LFInst_2_U7  ( .A(
        SubCellInst_LFInst_8_LFInst_2_n7 ), .B(AddKeyMUXOutput[34]), .Z(
        SubCellInst_LFInst_8_LFInst_2_n1 ) );
  ORN2 SubCellInst_LFInst_8_LFInst_2_U6  ( .A(AddKeyMUXOutput[33]), .B(
        AddKeyMUXOutput[35]), .Z(SubCellInst_LFInst_8_LFInst_2_n4 ) );
  AND2 SubCellInst_LFInst_8_LFInst_2_U5  ( .A(AddKeyMUXOutput[33]), .B(
        AddKeyMUXOutput[32]), .Z(SubCellInst_LFInst_8_LFInst_2_n6 ) );
  ORN2 SubCellInst_LFInst_8_LFInst_2_U4  ( .A(AddKeyMUXOutput[35]), .B(
        SubCellInst_LFInst_8_LFInst_2_n6 ), .Z(
        SubCellInst_LFInst_8_LFInst_2_n5 ) );
  AND2 SubCellInst_LFInst_8_LFInst_2_U3  ( .A(
        SubCellInst_LFInst_8_LFInst_2_n4 ), .B(
        SubCellInst_LFInst_8_LFInst_2_n5 ), .Z(
        SubCellInst_LFInst_8_LFInst_2_n3 ) );
  ORN2 SubCellInst_LFInst_8_LFInst_2_U2  ( .A(
        SubCellInst_LFInst_8_LFInst_2_n3 ), .B(AddKeyMUXOutput[34]), .Z(
        SubCellInst_LFInst_8_LFInst_2_n2 ) );
  ORN2 SubCellInst_LFInst_8_LFInst_2_U1  ( .A(
        SubCellInst_LFInst_8_LFInst_2_n1 ), .B(
        SubCellInst_LFInst_8_LFInst_2_n2 ), .Z(MCInst1_MC2_v1_3 [3]) );
  AND2 SubCellInst_LFInst_8_LFInst_1_U8  ( .A(AddKeyMUXOutput[34]), .B(
        AddKeyMUXOutput[32]), .Z(SubCellInst_LFInst_8_LFInst_1_n4 ) );
  AND2 SubCellInst_LFInst_8_LFInst_1_U7  ( .A(AddKeyMUXOutput[33]), .B(
        AddKeyMUXOutput[32]), .Z(SubCellInst_LFInst_8_LFInst_1_n7 ) );
  OR2 SubCellInst_LFInst_8_LFInst_1_U6  ( .A(AddKeyMUXOutput[34]), .B(
        SubCellInst_LFInst_8_LFInst_1_n7 ), .Z(
        SubCellInst_LFInst_8_LFInst_1_n6 ) );
  ORN2 SubCellInst_LFInst_8_LFInst_1_U5  ( .A(
        SubCellInst_LFInst_8_LFInst_1_n4 ), .B(
        SubCellInst_LFInst_8_LFInst_1_n6 ), .Z(
        SubCellInst_LFInst_8_LFInst_1_n5 ) );
  AND2 SubCellInst_LFInst_8_LFInst_1_U4  ( .A(AddKeyMUXOutput[35]), .B(
        SubCellInst_LFInst_8_LFInst_1_n5 ), .Z(
        SubCellInst_LFInst_8_LFInst_1_n1 ) );
  BIC2 SubCellInst_LFInst_8_LFInst_1_U3  ( .A(AddKeyMUXOutput[33]), .B(
        SubCellInst_LFInst_8_LFInst_1_n4 ), .Z(
        SubCellInst_LFInst_8_LFInst_1_n3 ) );
  ORN2 SubCellInst_LFInst_8_LFInst_1_U2  ( .A(AddKeyMUXOutput[35]), .B(
        SubCellInst_LFInst_8_LFInst_1_n3 ), .Z(
        SubCellInst_LFInst_8_LFInst_1_n2 ) );
  ORN2 SubCellInst_LFInst_8_LFInst_1_U1  ( .A(
        SubCellInst_LFInst_8_LFInst_1_n1 ), .B(
        SubCellInst_LFInst_8_LFInst_1_n2 ), .Z(MCInst1_MC2_v1_3 [2]) );
  BIC2 SubCellInst_LFInst_8_LFInst_0_U3  ( .A(AddKeyMUXOutput[34]), .B(
        AddKeyMUXOutput[33]), .Z(SubCellInst_LFInst_8_LFInst_0_n1 ) );
  XOR2 SubCellInst_LFInst_8_LFInst_0_U2  ( .A(AddKeyMUXOutput[35]), .B(
        AddKeyMUXOutput[32]), .Z(SubCellInst_LFInst_8_LFInst_0_n2 ) );
  XOR2 SubCellInst_LFInst_8_LFInst_0_U1  ( .A(
        SubCellInst_LFInst_8_LFInst_0_n1 ), .B(
        SubCellInst_LFInst_8_LFInst_0_n2 ), .Z(ShiftRowsOutput[36]) );
  OR2 SubCellInst_LFInst_9_LFInst_3_U9  ( .A(AddKeyMUXOutput[37]), .B(
        AddKeyMUXOutput[36]), .Z(SubCellInst_LFInst_9_LFInst_3_n5 ) );
  AND2 SubCellInst_LFInst_9_LFInst_3_U8  ( .A(AddKeyMUXOutput[39]), .B(
        SubCellInst_LFInst_9_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_9_LFInst_3_n7 ) );
  AND2 SubCellInst_LFInst_9_LFInst_3_U7  ( .A(AddKeyMUXOutput[36]), .B(
        AddKeyMUXOutput[37]), .Z(SubCellInst_LFInst_9_LFInst_3_n8 ) );
  OR2 SubCellInst_LFInst_9_LFInst_3_U6  ( .A(
        SubCellInst_LFInst_9_LFInst_3_n7 ), .B(
        SubCellInst_LFInst_9_LFInst_3_n8 ), .Z(
        SubCellInst_LFInst_9_LFInst_3_n6 ) );
  BIC2 SubCellInst_LFInst_9_LFInst_3_U5  ( .A(
        SubCellInst_LFInst_9_LFInst_3_n6 ), .B(AddKeyMUXOutput[38]), .Z(
        SubCellInst_LFInst_9_LFInst_3_n1 ) );
  AND2 SubCellInst_LFInst_9_LFInst_3_U4  ( .A(AddKeyMUXOutput[38]), .B(
        AddKeyMUXOutput[37]), .Z(SubCellInst_LFInst_9_LFInst_3_n4 ) );
  ORN2 SubCellInst_LFInst_9_LFInst_3_U3  ( .A(
        SubCellInst_LFInst_9_LFInst_3_n4 ), .B(
        SubCellInst_LFInst_9_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_9_LFInst_3_n3 ) );
  ORN2 SubCellInst_LFInst_9_LFInst_3_U2  ( .A(AddKeyMUXOutput[39]), .B(
        SubCellInst_LFInst_9_LFInst_3_n3 ), .Z(
        SubCellInst_LFInst_9_LFInst_3_n2 ) );
  ORN2 SubCellInst_LFInst_9_LFInst_3_U1  ( .A(
        SubCellInst_LFInst_9_LFInst_3_n1 ), .B(
        SubCellInst_LFInst_9_LFInst_3_n2 ), .Z(MCInst1_MC1_v1_3 [0]) );
  BIC2 SubCellInst_LFInst_9_LFInst_2_U11  ( .A(AddKeyMUXOutput[37]), .B(
        AddKeyMUXOutput[36]), .Z(SubCellInst_LFInst_9_LFInst_2_n8 ) );
  ORN2 SubCellInst_LFInst_9_LFInst_2_U10  ( .A(AddKeyMUXOutput[36]), .B(
        AddKeyMUXOutput[39]), .Z(SubCellInst_LFInst_9_LFInst_2_n10 ) );
  ORN2 SubCellInst_LFInst_9_LFInst_2_U9  ( .A(AddKeyMUXOutput[37]), .B(
        SubCellInst_LFInst_9_LFInst_2_n10 ), .Z(
        SubCellInst_LFInst_9_LFInst_2_n9 ) );
  ORN2 SubCellInst_LFInst_9_LFInst_2_U8  ( .A(
        SubCellInst_LFInst_9_LFInst_2_n8 ), .B(
        SubCellInst_LFInst_9_LFInst_2_n9 ), .Z(
        SubCellInst_LFInst_9_LFInst_2_n7 ) );
  BIC2 SubCellInst_LFInst_9_LFInst_2_U7  ( .A(
        SubCellInst_LFInst_9_LFInst_2_n7 ), .B(AddKeyMUXOutput[38]), .Z(
        SubCellInst_LFInst_9_LFInst_2_n1 ) );
  ORN2 SubCellInst_LFInst_9_LFInst_2_U6  ( .A(AddKeyMUXOutput[37]), .B(
        AddKeyMUXOutput[39]), .Z(SubCellInst_LFInst_9_LFInst_2_n4 ) );
  AND2 SubCellInst_LFInst_9_LFInst_2_U5  ( .A(AddKeyMUXOutput[37]), .B(
        AddKeyMUXOutput[36]), .Z(SubCellInst_LFInst_9_LFInst_2_n6 ) );
  ORN2 SubCellInst_LFInst_9_LFInst_2_U4  ( .A(AddKeyMUXOutput[39]), .B(
        SubCellInst_LFInst_9_LFInst_2_n6 ), .Z(
        SubCellInst_LFInst_9_LFInst_2_n5 ) );
  AND2 SubCellInst_LFInst_9_LFInst_2_U3  ( .A(
        SubCellInst_LFInst_9_LFInst_2_n4 ), .B(
        SubCellInst_LFInst_9_LFInst_2_n5 ), .Z(
        SubCellInst_LFInst_9_LFInst_2_n3 ) );
  ORN2 SubCellInst_LFInst_9_LFInst_2_U2  ( .A(
        SubCellInst_LFInst_9_LFInst_2_n3 ), .B(AddKeyMUXOutput[38]), .Z(
        SubCellInst_LFInst_9_LFInst_2_n2 ) );
  ORN2 SubCellInst_LFInst_9_LFInst_2_U1  ( .A(
        SubCellInst_LFInst_9_LFInst_2_n1 ), .B(
        SubCellInst_LFInst_9_LFInst_2_n2 ), .Z(MCInst1_MC1_v1_3 [3]) );
  AND2 SubCellInst_LFInst_9_LFInst_1_U8  ( .A(AddKeyMUXOutput[38]), .B(
        AddKeyMUXOutput[36]), .Z(SubCellInst_LFInst_9_LFInst_1_n4 ) );
  AND2 SubCellInst_LFInst_9_LFInst_1_U7  ( .A(AddKeyMUXOutput[37]), .B(
        AddKeyMUXOutput[36]), .Z(SubCellInst_LFInst_9_LFInst_1_n7 ) );
  OR2 SubCellInst_LFInst_9_LFInst_1_U6  ( .A(AddKeyMUXOutput[38]), .B(
        SubCellInst_LFInst_9_LFInst_1_n7 ), .Z(
        SubCellInst_LFInst_9_LFInst_1_n6 ) );
  ORN2 SubCellInst_LFInst_9_LFInst_1_U5  ( .A(
        SubCellInst_LFInst_9_LFInst_1_n4 ), .B(
        SubCellInst_LFInst_9_LFInst_1_n6 ), .Z(
        SubCellInst_LFInst_9_LFInst_1_n5 ) );
  AND2 SubCellInst_LFInst_9_LFInst_1_U4  ( .A(AddKeyMUXOutput[39]), .B(
        SubCellInst_LFInst_9_LFInst_1_n5 ), .Z(
        SubCellInst_LFInst_9_LFInst_1_n1 ) );
  BIC2 SubCellInst_LFInst_9_LFInst_1_U3  ( .A(AddKeyMUXOutput[37]), .B(
        SubCellInst_LFInst_9_LFInst_1_n4 ), .Z(
        SubCellInst_LFInst_9_LFInst_1_n3 ) );
  ORN2 SubCellInst_LFInst_9_LFInst_1_U2  ( .A(AddKeyMUXOutput[39]), .B(
        SubCellInst_LFInst_9_LFInst_1_n3 ), .Z(
        SubCellInst_LFInst_9_LFInst_1_n2 ) );
  ORN2 SubCellInst_LFInst_9_LFInst_1_U1  ( .A(
        SubCellInst_LFInst_9_LFInst_1_n1 ), .B(
        SubCellInst_LFInst_9_LFInst_1_n2 ), .Z(MCInst1_MC1_v1_3 [2]) );
  BIC2 SubCellInst_LFInst_9_LFInst_0_U3  ( .A(AddKeyMUXOutput[38]), .B(
        AddKeyMUXOutput[37]), .Z(SubCellInst_LFInst_9_LFInst_0_n1 ) );
  XOR2 SubCellInst_LFInst_9_LFInst_0_U2  ( .A(AddKeyMUXOutput[39]), .B(
        AddKeyMUXOutput[36]), .Z(SubCellInst_LFInst_9_LFInst_0_n2 ) );
  XOR2 SubCellInst_LFInst_9_LFInst_0_U1  ( .A(
        SubCellInst_LFInst_9_LFInst_0_n1 ), .B(
        SubCellInst_LFInst_9_LFInst_0_n2 ), .Z(ShiftRowsOutput[40]) );
  OR2 SubCellInst_LFInst_10_LFInst_3_U9  ( .A(AddConstOutput[17]), .B(
        AddConstOutput[16]), .Z(SubCellInst_LFInst_10_LFInst_3_n5 ) );
  AND2 SubCellInst_LFInst_10_LFInst_3_U8  ( .A(AddConstOutput[19]), .B(
        SubCellInst_LFInst_10_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_10_LFInst_3_n7 ) );
  AND2 SubCellInst_LFInst_10_LFInst_3_U7  ( .A(AddConstOutput[16]), .B(
        AddConstOutput[17]), .Z(SubCellInst_LFInst_10_LFInst_3_n8 ) );
  OR2 SubCellInst_LFInst_10_LFInst_3_U6  ( .A(
        SubCellInst_LFInst_10_LFInst_3_n7 ), .B(
        SubCellInst_LFInst_10_LFInst_3_n8 ), .Z(
        SubCellInst_LFInst_10_LFInst_3_n6 ) );
  BIC2 SubCellInst_LFInst_10_LFInst_3_U5  ( .A(
        SubCellInst_LFInst_10_LFInst_3_n6 ), .B(AddConstOutput[18]), .Z(
        SubCellInst_LFInst_10_LFInst_3_n1 ) );
  AND2 SubCellInst_LFInst_10_LFInst_3_U4  ( .A(AddConstOutput[18]), .B(
        AddConstOutput[17]), .Z(SubCellInst_LFInst_10_LFInst_3_n4 ) );
  ORN2 SubCellInst_LFInst_10_LFInst_3_U3  ( .A(
        SubCellInst_LFInst_10_LFInst_3_n4 ), .B(
        SubCellInst_LFInst_10_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_10_LFInst_3_n3 ) );
  ORN2 SubCellInst_LFInst_10_LFInst_3_U2  ( .A(AddConstOutput[19]), .B(
        SubCellInst_LFInst_10_LFInst_3_n3 ), .Z(
        SubCellInst_LFInst_10_LFInst_3_n2 ) );
  ORN2 SubCellInst_LFInst_10_LFInst_3_U1  ( .A(
        SubCellInst_LFInst_10_LFInst_3_n1 ), .B(
        SubCellInst_LFInst_10_LFInst_3_n2 ), .Z(MCInst1_MC0_v1_3 [0]) );
  BIC2 SubCellInst_LFInst_10_LFInst_2_U11  ( .A(AddConstOutput[17]), .B(
        AddConstOutput[16]), .Z(SubCellInst_LFInst_10_LFInst_2_n8 ) );
  ORN2 SubCellInst_LFInst_10_LFInst_2_U10  ( .A(AddConstOutput[16]), .B(
        AddConstOutput[19]), .Z(SubCellInst_LFInst_10_LFInst_2_n10 ) );
  ORN2 SubCellInst_LFInst_10_LFInst_2_U9  ( .A(AddConstOutput[17]), .B(
        SubCellInst_LFInst_10_LFInst_2_n10 ), .Z(
        SubCellInst_LFInst_10_LFInst_2_n9 ) );
  ORN2 SubCellInst_LFInst_10_LFInst_2_U8  ( .A(
        SubCellInst_LFInst_10_LFInst_2_n8 ), .B(
        SubCellInst_LFInst_10_LFInst_2_n9 ), .Z(
        SubCellInst_LFInst_10_LFInst_2_n7 ) );
  BIC2 SubCellInst_LFInst_10_LFInst_2_U7  ( .A(
        SubCellInst_LFInst_10_LFInst_2_n7 ), .B(AddConstOutput[18]), .Z(
        SubCellInst_LFInst_10_LFInst_2_n1 ) );
  ORN2 SubCellInst_LFInst_10_LFInst_2_U6  ( .A(AddConstOutput[17]), .B(
        AddConstOutput[19]), .Z(SubCellInst_LFInst_10_LFInst_2_n4 ) );
  AND2 SubCellInst_LFInst_10_LFInst_2_U5  ( .A(AddConstOutput[17]), .B(
        AddConstOutput[16]), .Z(SubCellInst_LFInst_10_LFInst_2_n6 ) );
  ORN2 SubCellInst_LFInst_10_LFInst_2_U4  ( .A(AddConstOutput[19]), .B(
        SubCellInst_LFInst_10_LFInst_2_n6 ), .Z(
        SubCellInst_LFInst_10_LFInst_2_n5 ) );
  AND2 SubCellInst_LFInst_10_LFInst_2_U3  ( .A(
        SubCellInst_LFInst_10_LFInst_2_n4 ), .B(
        SubCellInst_LFInst_10_LFInst_2_n5 ), .Z(
        SubCellInst_LFInst_10_LFInst_2_n3 ) );
  ORN2 SubCellInst_LFInst_10_LFInst_2_U2  ( .A(
        SubCellInst_LFInst_10_LFInst_2_n3 ), .B(AddConstOutput[18]), .Z(
        SubCellInst_LFInst_10_LFInst_2_n2 ) );
  ORN2 SubCellInst_LFInst_10_LFInst_2_U1  ( .A(
        SubCellInst_LFInst_10_LFInst_2_n1 ), .B(
        SubCellInst_LFInst_10_LFInst_2_n2 ), .Z(MCInst1_MC0_v1_3 [3]) );
  AND2 SubCellInst_LFInst_10_LFInst_1_U8  ( .A(AddConstOutput[18]), .B(
        AddConstOutput[16]), .Z(SubCellInst_LFInst_10_LFInst_1_n4 ) );
  AND2 SubCellInst_LFInst_10_LFInst_1_U7  ( .A(AddConstOutput[17]), .B(
        AddConstOutput[16]), .Z(SubCellInst_LFInst_10_LFInst_1_n7 ) );
  OR2 SubCellInst_LFInst_10_LFInst_1_U6  ( .A(AddConstOutput[18]), .B(
        SubCellInst_LFInst_10_LFInst_1_n7 ), .Z(
        SubCellInst_LFInst_10_LFInst_1_n6 ) );
  ORN2 SubCellInst_LFInst_10_LFInst_1_U5  ( .A(
        SubCellInst_LFInst_10_LFInst_1_n4 ), .B(
        SubCellInst_LFInst_10_LFInst_1_n6 ), .Z(
        SubCellInst_LFInst_10_LFInst_1_n5 ) );
  AND2 SubCellInst_LFInst_10_LFInst_1_U4  ( .A(AddConstOutput[19]), .B(
        SubCellInst_LFInst_10_LFInst_1_n5 ), .Z(
        SubCellInst_LFInst_10_LFInst_1_n1 ) );
  BIC2 SubCellInst_LFInst_10_LFInst_1_U3  ( .A(AddConstOutput[17]), .B(
        SubCellInst_LFInst_10_LFInst_1_n4 ), .Z(
        SubCellInst_LFInst_10_LFInst_1_n3 ) );
  ORN2 SubCellInst_LFInst_10_LFInst_1_U2  ( .A(AddConstOutput[19]), .B(
        SubCellInst_LFInst_10_LFInst_1_n3 ), .Z(
        SubCellInst_LFInst_10_LFInst_1_n2 ) );
  ORN2 SubCellInst_LFInst_10_LFInst_1_U1  ( .A(
        SubCellInst_LFInst_10_LFInst_1_n1 ), .B(
        SubCellInst_LFInst_10_LFInst_1_n2 ), .Z(MCInst1_MC0_v1_3 [2]) );
  BIC2 SubCellInst_LFInst_10_LFInst_0_U3  ( .A(AddConstOutput[18]), .B(
        AddConstOutput[17]), .Z(SubCellInst_LFInst_10_LFInst_0_n1 ) );
  XOR2 SubCellInst_LFInst_10_LFInst_0_U2  ( .A(AddConstOutput[19]), .B(
        AddConstOutput[16]), .Z(SubCellInst_LFInst_10_LFInst_0_n2 ) );
  XOR2 SubCellInst_LFInst_10_LFInst_0_U1  ( .A(
        SubCellInst_LFInst_10_LFInst_0_n1 ), .B(
        SubCellInst_LFInst_10_LFInst_0_n2 ), .Z(ShiftRowsOutput[44]) );
  OR2 SubCellInst_LFInst_11_LFInst_3_U9  ( .A(AddConstOutput[21]), .B(
        AddConstOutput[20]), .Z(SubCellInst_LFInst_11_LFInst_3_n5 ) );
  AND2 SubCellInst_LFInst_11_LFInst_3_U8  ( .A(AddConstOutput[23]), .B(
        SubCellInst_LFInst_11_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_11_LFInst_3_n7 ) );
  AND2 SubCellInst_LFInst_11_LFInst_3_U7  ( .A(AddConstOutput[20]), .B(
        AddConstOutput[21]), .Z(SubCellInst_LFInst_11_LFInst_3_n8 ) );
  OR2 SubCellInst_LFInst_11_LFInst_3_U6  ( .A(
        SubCellInst_LFInst_11_LFInst_3_n7 ), .B(
        SubCellInst_LFInst_11_LFInst_3_n8 ), .Z(
        SubCellInst_LFInst_11_LFInst_3_n6 ) );
  BIC2 SubCellInst_LFInst_11_LFInst_3_U5  ( .A(
        SubCellInst_LFInst_11_LFInst_3_n6 ), .B(AddConstOutput[22]), .Z(
        SubCellInst_LFInst_11_LFInst_3_n1 ) );
  AND2 SubCellInst_LFInst_11_LFInst_3_U4  ( .A(AddConstOutput[22]), .B(
        AddConstOutput[21]), .Z(SubCellInst_LFInst_11_LFInst_3_n4 ) );
  ORN2 SubCellInst_LFInst_11_LFInst_3_U3  ( .A(
        SubCellInst_LFInst_11_LFInst_3_n4 ), .B(
        SubCellInst_LFInst_11_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_11_LFInst_3_n3 ) );
  ORN2 SubCellInst_LFInst_11_LFInst_3_U2  ( .A(AddConstOutput[23]), .B(
        SubCellInst_LFInst_11_LFInst_3_n3 ), .Z(
        SubCellInst_LFInst_11_LFInst_3_n2 ) );
  ORN2 SubCellInst_LFInst_11_LFInst_3_U1  ( .A(
        SubCellInst_LFInst_11_LFInst_3_n1 ), .B(
        SubCellInst_LFInst_11_LFInst_3_n2 ), .Z(MCInst1_MC3_v1_3 [0]) );
  BIC2 SubCellInst_LFInst_11_LFInst_2_U11  ( .A(AddConstOutput[21]), .B(
        AddConstOutput[20]), .Z(SubCellInst_LFInst_11_LFInst_2_n8 ) );
  ORN2 SubCellInst_LFInst_11_LFInst_2_U10  ( .A(AddConstOutput[20]), .B(
        AddConstOutput[23]), .Z(SubCellInst_LFInst_11_LFInst_2_n10 ) );
  ORN2 SubCellInst_LFInst_11_LFInst_2_U9  ( .A(AddConstOutput[21]), .B(
        SubCellInst_LFInst_11_LFInst_2_n10 ), .Z(
        SubCellInst_LFInst_11_LFInst_2_n9 ) );
  ORN2 SubCellInst_LFInst_11_LFInst_2_U8  ( .A(
        SubCellInst_LFInst_11_LFInst_2_n8 ), .B(
        SubCellInst_LFInst_11_LFInst_2_n9 ), .Z(
        SubCellInst_LFInst_11_LFInst_2_n7 ) );
  BIC2 SubCellInst_LFInst_11_LFInst_2_U7  ( .A(
        SubCellInst_LFInst_11_LFInst_2_n7 ), .B(AddConstOutput[22]), .Z(
        SubCellInst_LFInst_11_LFInst_2_n1 ) );
  ORN2 SubCellInst_LFInst_11_LFInst_2_U6  ( .A(AddConstOutput[21]), .B(
        AddConstOutput[23]), .Z(SubCellInst_LFInst_11_LFInst_2_n4 ) );
  AND2 SubCellInst_LFInst_11_LFInst_2_U5  ( .A(AddConstOutput[21]), .B(
        AddConstOutput[20]), .Z(SubCellInst_LFInst_11_LFInst_2_n6 ) );
  ORN2 SubCellInst_LFInst_11_LFInst_2_U4  ( .A(AddConstOutput[23]), .B(
        SubCellInst_LFInst_11_LFInst_2_n6 ), .Z(
        SubCellInst_LFInst_11_LFInst_2_n5 ) );
  AND2 SubCellInst_LFInst_11_LFInst_2_U3  ( .A(
        SubCellInst_LFInst_11_LFInst_2_n4 ), .B(
        SubCellInst_LFInst_11_LFInst_2_n5 ), .Z(
        SubCellInst_LFInst_11_LFInst_2_n3 ) );
  ORN2 SubCellInst_LFInst_11_LFInst_2_U2  ( .A(
        SubCellInst_LFInst_11_LFInst_2_n3 ), .B(AddConstOutput[22]), .Z(
        SubCellInst_LFInst_11_LFInst_2_n2 ) );
  ORN2 SubCellInst_LFInst_11_LFInst_2_U1  ( .A(
        SubCellInst_LFInst_11_LFInst_2_n1 ), .B(
        SubCellInst_LFInst_11_LFInst_2_n2 ), .Z(MCInst1_MC3_v1_3 [3]) );
  AND2 SubCellInst_LFInst_11_LFInst_1_U8  ( .A(AddConstOutput[22]), .B(
        AddConstOutput[20]), .Z(SubCellInst_LFInst_11_LFInst_1_n4 ) );
  AND2 SubCellInst_LFInst_11_LFInst_1_U7  ( .A(AddConstOutput[21]), .B(
        AddConstOutput[20]), .Z(SubCellInst_LFInst_11_LFInst_1_n7 ) );
  OR2 SubCellInst_LFInst_11_LFInst_1_U6  ( .A(AddConstOutput[22]), .B(
        SubCellInst_LFInst_11_LFInst_1_n7 ), .Z(
        SubCellInst_LFInst_11_LFInst_1_n6 ) );
  ORN2 SubCellInst_LFInst_11_LFInst_1_U5  ( .A(
        SubCellInst_LFInst_11_LFInst_1_n4 ), .B(
        SubCellInst_LFInst_11_LFInst_1_n6 ), .Z(
        SubCellInst_LFInst_11_LFInst_1_n5 ) );
  AND2 SubCellInst_LFInst_11_LFInst_1_U4  ( .A(AddConstOutput[23]), .B(
        SubCellInst_LFInst_11_LFInst_1_n5 ), .Z(
        SubCellInst_LFInst_11_LFInst_1_n1 ) );
  BIC2 SubCellInst_LFInst_11_LFInst_1_U3  ( .A(AddConstOutput[21]), .B(
        SubCellInst_LFInst_11_LFInst_1_n4 ), .Z(
        SubCellInst_LFInst_11_LFInst_1_n3 ) );
  ORN2 SubCellInst_LFInst_11_LFInst_1_U2  ( .A(AddConstOutput[23]), .B(
        SubCellInst_LFInst_11_LFInst_1_n3 ), .Z(
        SubCellInst_LFInst_11_LFInst_1_n2 ) );
  ORN2 SubCellInst_LFInst_11_LFInst_1_U1  ( .A(
        SubCellInst_LFInst_11_LFInst_1_n1 ), .B(
        SubCellInst_LFInst_11_LFInst_1_n2 ), .Z(MCInst1_MC3_v1_3 [2]) );
  BIC2 SubCellInst_LFInst_11_LFInst_0_U3  ( .A(AddConstOutput[22]), .B(
        AddConstOutput[21]), .Z(SubCellInst_LFInst_11_LFInst_0_n1 ) );
  XOR2 SubCellInst_LFInst_11_LFInst_0_U2  ( .A(AddConstOutput[23]), .B(
        AddConstOutput[20]), .Z(SubCellInst_LFInst_11_LFInst_0_n2 ) );
  XOR2 SubCellInst_LFInst_11_LFInst_0_U1  ( .A(
        SubCellInst_LFInst_11_LFInst_0_n1 ), .B(
        SubCellInst_LFInst_11_LFInst_0_n2 ), .Z(ShiftRowsOutput[32]) );
  OR2 SubCellInst_LFInst_12_LFInst_3_U9  ( .A(AddKeyMUXOutput[49]), .B(
        AddKeyMUXOutput[48]), .Z(SubCellInst_LFInst_12_LFInst_3_n5 ) );
  AND2 SubCellInst_LFInst_12_LFInst_3_U8  ( .A(AddKeyMUXOutput[51]), .B(
        SubCellInst_LFInst_12_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_12_LFInst_3_n7 ) );
  AND2 SubCellInst_LFInst_12_LFInst_3_U7  ( .A(AddKeyMUXOutput[48]), .B(
        AddKeyMUXOutput[49]), .Z(SubCellInst_LFInst_12_LFInst_3_n8 ) );
  OR2 SubCellInst_LFInst_12_LFInst_3_U6  ( .A(
        SubCellInst_LFInst_12_LFInst_3_n7 ), .B(
        SubCellInst_LFInst_12_LFInst_3_n8 ), .Z(
        SubCellInst_LFInst_12_LFInst_3_n6 ) );
  BIC2 SubCellInst_LFInst_12_LFInst_3_U5  ( .A(
        SubCellInst_LFInst_12_LFInst_3_n6 ), .B(AddKeyMUXOutput[50]), .Z(
        SubCellInst_LFInst_12_LFInst_3_n1 ) );
  AND2 SubCellInst_LFInst_12_LFInst_3_U4  ( .A(AddKeyMUXOutput[50]), .B(
        AddKeyMUXOutput[49]), .Z(SubCellInst_LFInst_12_LFInst_3_n4 ) );
  ORN2 SubCellInst_LFInst_12_LFInst_3_U3  ( .A(
        SubCellInst_LFInst_12_LFInst_3_n4 ), .B(
        SubCellInst_LFInst_12_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_12_LFInst_3_n3 ) );
  ORN2 SubCellInst_LFInst_12_LFInst_3_U2  ( .A(AddKeyMUXOutput[51]), .B(
        SubCellInst_LFInst_12_LFInst_3_n3 ), .Z(
        SubCellInst_LFInst_12_LFInst_3_n2 ) );
  ORN2 SubCellInst_LFInst_12_LFInst_3_U1  ( .A(
        SubCellInst_LFInst_12_LFInst_3_n1 ), .B(
        SubCellInst_LFInst_12_LFInst_3_n2 ), .Z(MCInst1_MC3_v0_3 [0]) );
  BIC2 SubCellInst_LFInst_12_LFInst_2_U11  ( .A(AddKeyMUXOutput[49]), .B(
        AddKeyMUXOutput[48]), .Z(SubCellInst_LFInst_12_LFInst_2_n8 ) );
  ORN2 SubCellInst_LFInst_12_LFInst_2_U10  ( .A(AddKeyMUXOutput[48]), .B(
        AddKeyMUXOutput[51]), .Z(SubCellInst_LFInst_12_LFInst_2_n10 ) );
  ORN2 SubCellInst_LFInst_12_LFInst_2_U9  ( .A(AddKeyMUXOutput[49]), .B(
        SubCellInst_LFInst_12_LFInst_2_n10 ), .Z(
        SubCellInst_LFInst_12_LFInst_2_n9 ) );
  ORN2 SubCellInst_LFInst_12_LFInst_2_U8  ( .A(
        SubCellInst_LFInst_12_LFInst_2_n8 ), .B(
        SubCellInst_LFInst_12_LFInst_2_n9 ), .Z(
        SubCellInst_LFInst_12_LFInst_2_n7 ) );
  BIC2 SubCellInst_LFInst_12_LFInst_2_U7  ( .A(
        SubCellInst_LFInst_12_LFInst_2_n7 ), .B(AddKeyMUXOutput[50]), .Z(
        SubCellInst_LFInst_12_LFInst_2_n1 ) );
  ORN2 SubCellInst_LFInst_12_LFInst_2_U6  ( .A(AddKeyMUXOutput[49]), .B(
        AddKeyMUXOutput[51]), .Z(SubCellInst_LFInst_12_LFInst_2_n4 ) );
  AND2 SubCellInst_LFInst_12_LFInst_2_U5  ( .A(AddKeyMUXOutput[49]), .B(
        AddKeyMUXOutput[48]), .Z(SubCellInst_LFInst_12_LFInst_2_n6 ) );
  ORN2 SubCellInst_LFInst_12_LFInst_2_U4  ( .A(AddKeyMUXOutput[51]), .B(
        SubCellInst_LFInst_12_LFInst_2_n6 ), .Z(
        SubCellInst_LFInst_12_LFInst_2_n5 ) );
  AND2 SubCellInst_LFInst_12_LFInst_2_U3  ( .A(
        SubCellInst_LFInst_12_LFInst_2_n4 ), .B(
        SubCellInst_LFInst_12_LFInst_2_n5 ), .Z(
        SubCellInst_LFInst_12_LFInst_2_n3 ) );
  ORN2 SubCellInst_LFInst_12_LFInst_2_U2  ( .A(
        SubCellInst_LFInst_12_LFInst_2_n3 ), .B(AddKeyMUXOutput[50]), .Z(
        SubCellInst_LFInst_12_LFInst_2_n2 ) );
  ORN2 SubCellInst_LFInst_12_LFInst_2_U1  ( .A(
        SubCellInst_LFInst_12_LFInst_2_n1 ), .B(
        SubCellInst_LFInst_12_LFInst_2_n2 ), .Z(MCInst1_MC3_v0_3 [3]) );
  AND2 SubCellInst_LFInst_12_LFInst_1_U8  ( .A(AddKeyMUXOutput[50]), .B(
        AddKeyMUXOutput[48]), .Z(SubCellInst_LFInst_12_LFInst_1_n4 ) );
  AND2 SubCellInst_LFInst_12_LFInst_1_U7  ( .A(AddKeyMUXOutput[49]), .B(
        AddKeyMUXOutput[48]), .Z(SubCellInst_LFInst_12_LFInst_1_n7 ) );
  OR2 SubCellInst_LFInst_12_LFInst_1_U6  ( .A(AddKeyMUXOutput[50]), .B(
        SubCellInst_LFInst_12_LFInst_1_n7 ), .Z(
        SubCellInst_LFInst_12_LFInst_1_n6 ) );
  ORN2 SubCellInst_LFInst_12_LFInst_1_U5  ( .A(
        SubCellInst_LFInst_12_LFInst_1_n4 ), .B(
        SubCellInst_LFInst_12_LFInst_1_n6 ), .Z(
        SubCellInst_LFInst_12_LFInst_1_n5 ) );
  AND2 SubCellInst_LFInst_12_LFInst_1_U4  ( .A(AddKeyMUXOutput[51]), .B(
        SubCellInst_LFInst_12_LFInst_1_n5 ), .Z(
        SubCellInst_LFInst_12_LFInst_1_n1 ) );
  BIC2 SubCellInst_LFInst_12_LFInst_1_U3  ( .A(AddKeyMUXOutput[49]), .B(
        SubCellInst_LFInst_12_LFInst_1_n4 ), .Z(
        SubCellInst_LFInst_12_LFInst_1_n3 ) );
  ORN2 SubCellInst_LFInst_12_LFInst_1_U2  ( .A(AddKeyMUXOutput[51]), .B(
        SubCellInst_LFInst_12_LFInst_1_n3 ), .Z(
        SubCellInst_LFInst_12_LFInst_1_n2 ) );
  ORN2 SubCellInst_LFInst_12_LFInst_1_U1  ( .A(
        SubCellInst_LFInst_12_LFInst_1_n1 ), .B(
        SubCellInst_LFInst_12_LFInst_1_n2 ), .Z(MCInst1_MC3_v0_0 [3]) );
  BIC2 SubCellInst_LFInst_12_LFInst_0_U3  ( .A(AddKeyMUXOutput[50]), .B(
        AddKeyMUXOutput[49]), .Z(SubCellInst_LFInst_12_LFInst_0_n1 ) );
  XOR2 SubCellInst_LFInst_12_LFInst_0_U2  ( .A(AddKeyMUXOutput[51]), .B(
        AddKeyMUXOutput[48]), .Z(SubCellInst_LFInst_12_LFInst_0_n2 ) );
  XOR2 SubCellInst_LFInst_12_LFInst_0_U1  ( .A(
        SubCellInst_LFInst_12_LFInst_0_n1 ), .B(
        SubCellInst_LFInst_12_LFInst_0_n2 ), .Z(ShiftRowsOutput[48]) );
  OR2 SubCellInst_LFInst_13_LFInst_3_U9  ( .A(AddKeyMUXOutput[53]), .B(
        AddKeyMUXOutput[52]), .Z(SubCellInst_LFInst_13_LFInst_3_n5 ) );
  AND2 SubCellInst_LFInst_13_LFInst_3_U8  ( .A(AddKeyMUXOutput[55]), .B(
        SubCellInst_LFInst_13_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_13_LFInst_3_n7 ) );
  AND2 SubCellInst_LFInst_13_LFInst_3_U7  ( .A(AddKeyMUXOutput[52]), .B(
        AddKeyMUXOutput[53]), .Z(SubCellInst_LFInst_13_LFInst_3_n8 ) );
  OR2 SubCellInst_LFInst_13_LFInst_3_U6  ( .A(
        SubCellInst_LFInst_13_LFInst_3_n7 ), .B(
        SubCellInst_LFInst_13_LFInst_3_n8 ), .Z(
        SubCellInst_LFInst_13_LFInst_3_n6 ) );
  BIC2 SubCellInst_LFInst_13_LFInst_3_U5  ( .A(
        SubCellInst_LFInst_13_LFInst_3_n6 ), .B(AddKeyMUXOutput[54]), .Z(
        SubCellInst_LFInst_13_LFInst_3_n1 ) );
  AND2 SubCellInst_LFInst_13_LFInst_3_U4  ( .A(AddKeyMUXOutput[54]), .B(
        AddKeyMUXOutput[53]), .Z(SubCellInst_LFInst_13_LFInst_3_n4 ) );
  ORN2 SubCellInst_LFInst_13_LFInst_3_U3  ( .A(
        SubCellInst_LFInst_13_LFInst_3_n4 ), .B(
        SubCellInst_LFInst_13_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_13_LFInst_3_n3 ) );
  ORN2 SubCellInst_LFInst_13_LFInst_3_U2  ( .A(AddKeyMUXOutput[55]), .B(
        SubCellInst_LFInst_13_LFInst_3_n3 ), .Z(
        SubCellInst_LFInst_13_LFInst_3_n2 ) );
  ORN2 SubCellInst_LFInst_13_LFInst_3_U1  ( .A(
        SubCellInst_LFInst_13_LFInst_3_n1 ), .B(
        SubCellInst_LFInst_13_LFInst_3_n2 ), .Z(MCInst1_MC2_v0_3 [0]) );
  BIC2 SubCellInst_LFInst_13_LFInst_2_U11  ( .A(AddKeyMUXOutput[53]), .B(
        AddKeyMUXOutput[52]), .Z(SubCellInst_LFInst_13_LFInst_2_n8 ) );
  ORN2 SubCellInst_LFInst_13_LFInst_2_U10  ( .A(AddKeyMUXOutput[52]), .B(
        AddKeyMUXOutput[55]), .Z(SubCellInst_LFInst_13_LFInst_2_n10 ) );
  ORN2 SubCellInst_LFInst_13_LFInst_2_U9  ( .A(AddKeyMUXOutput[53]), .B(
        SubCellInst_LFInst_13_LFInst_2_n10 ), .Z(
        SubCellInst_LFInst_13_LFInst_2_n9 ) );
  ORN2 SubCellInst_LFInst_13_LFInst_2_U8  ( .A(
        SubCellInst_LFInst_13_LFInst_2_n8 ), .B(
        SubCellInst_LFInst_13_LFInst_2_n9 ), .Z(
        SubCellInst_LFInst_13_LFInst_2_n7 ) );
  BIC2 SubCellInst_LFInst_13_LFInst_2_U7  ( .A(
        SubCellInst_LFInst_13_LFInst_2_n7 ), .B(AddKeyMUXOutput[54]), .Z(
        SubCellInst_LFInst_13_LFInst_2_n1 ) );
  ORN2 SubCellInst_LFInst_13_LFInst_2_U6  ( .A(AddKeyMUXOutput[53]), .B(
        AddKeyMUXOutput[55]), .Z(SubCellInst_LFInst_13_LFInst_2_n4 ) );
  AND2 SubCellInst_LFInst_13_LFInst_2_U5  ( .A(AddKeyMUXOutput[53]), .B(
        AddKeyMUXOutput[52]), .Z(SubCellInst_LFInst_13_LFInst_2_n6 ) );
  ORN2 SubCellInst_LFInst_13_LFInst_2_U4  ( .A(AddKeyMUXOutput[55]), .B(
        SubCellInst_LFInst_13_LFInst_2_n6 ), .Z(
        SubCellInst_LFInst_13_LFInst_2_n5 ) );
  AND2 SubCellInst_LFInst_13_LFInst_2_U3  ( .A(
        SubCellInst_LFInst_13_LFInst_2_n4 ), .B(
        SubCellInst_LFInst_13_LFInst_2_n5 ), .Z(
        SubCellInst_LFInst_13_LFInst_2_n3 ) );
  ORN2 SubCellInst_LFInst_13_LFInst_2_U2  ( .A(
        SubCellInst_LFInst_13_LFInst_2_n3 ), .B(AddKeyMUXOutput[54]), .Z(
        SubCellInst_LFInst_13_LFInst_2_n2 ) );
  ORN2 SubCellInst_LFInst_13_LFInst_2_U1  ( .A(
        SubCellInst_LFInst_13_LFInst_2_n1 ), .B(
        SubCellInst_LFInst_13_LFInst_2_n2 ), .Z(MCInst1_MC2_v0_3 [3]) );
  AND2 SubCellInst_LFInst_13_LFInst_1_U8  ( .A(AddKeyMUXOutput[54]), .B(
        AddKeyMUXOutput[52]), .Z(SubCellInst_LFInst_13_LFInst_1_n4 ) );
  AND2 SubCellInst_LFInst_13_LFInst_1_U7  ( .A(AddKeyMUXOutput[53]), .B(
        AddKeyMUXOutput[52]), .Z(SubCellInst_LFInst_13_LFInst_1_n7 ) );
  OR2 SubCellInst_LFInst_13_LFInst_1_U6  ( .A(AddKeyMUXOutput[54]), .B(
        SubCellInst_LFInst_13_LFInst_1_n7 ), .Z(
        SubCellInst_LFInst_13_LFInst_1_n6 ) );
  ORN2 SubCellInst_LFInst_13_LFInst_1_U5  ( .A(
        SubCellInst_LFInst_13_LFInst_1_n4 ), .B(
        SubCellInst_LFInst_13_LFInst_1_n6 ), .Z(
        SubCellInst_LFInst_13_LFInst_1_n5 ) );
  AND2 SubCellInst_LFInst_13_LFInst_1_U4  ( .A(AddKeyMUXOutput[55]), .B(
        SubCellInst_LFInst_13_LFInst_1_n5 ), .Z(
        SubCellInst_LFInst_13_LFInst_1_n1 ) );
  BIC2 SubCellInst_LFInst_13_LFInst_1_U3  ( .A(AddKeyMUXOutput[53]), .B(
        SubCellInst_LFInst_13_LFInst_1_n4 ), .Z(
        SubCellInst_LFInst_13_LFInst_1_n3 ) );
  ORN2 SubCellInst_LFInst_13_LFInst_1_U2  ( .A(AddKeyMUXOutput[55]), .B(
        SubCellInst_LFInst_13_LFInst_1_n3 ), .Z(
        SubCellInst_LFInst_13_LFInst_1_n2 ) );
  ORN2 SubCellInst_LFInst_13_LFInst_1_U1  ( .A(
        SubCellInst_LFInst_13_LFInst_1_n1 ), .B(
        SubCellInst_LFInst_13_LFInst_1_n2 ), .Z(MCInst1_MC2_v0_0 [3]) );
  BIC2 SubCellInst_LFInst_13_LFInst_0_U3  ( .A(AddKeyMUXOutput[54]), .B(
        AddKeyMUXOutput[53]), .Z(SubCellInst_LFInst_13_LFInst_0_n1 ) );
  XOR2 SubCellInst_LFInst_13_LFInst_0_U2  ( .A(AddKeyMUXOutput[55]), .B(
        AddKeyMUXOutput[52]), .Z(SubCellInst_LFInst_13_LFInst_0_n2 ) );
  XOR2 SubCellInst_LFInst_13_LFInst_0_U1  ( .A(
        SubCellInst_LFInst_13_LFInst_0_n1 ), .B(
        SubCellInst_LFInst_13_LFInst_0_n2 ), .Z(ShiftRowsOutput[52]) );
  OR2 SubCellInst_LFInst_14_LFInst_3_U9  ( .A(AddConstOutput[25]), .B(
        AddConstOutput[24]), .Z(SubCellInst_LFInst_14_LFInst_3_n5 ) );
  AND2 SubCellInst_LFInst_14_LFInst_3_U8  ( .A(AddConstOutput[27]), .B(
        SubCellInst_LFInst_14_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_14_LFInst_3_n7 ) );
  AND2 SubCellInst_LFInst_14_LFInst_3_U7  ( .A(AddConstOutput[24]), .B(
        AddConstOutput[25]), .Z(SubCellInst_LFInst_14_LFInst_3_n8 ) );
  OR2 SubCellInst_LFInst_14_LFInst_3_U6  ( .A(
        SubCellInst_LFInst_14_LFInst_3_n7 ), .B(
        SubCellInst_LFInst_14_LFInst_3_n8 ), .Z(
        SubCellInst_LFInst_14_LFInst_3_n6 ) );
  BIC2 SubCellInst_LFInst_14_LFInst_3_U5  ( .A(
        SubCellInst_LFInst_14_LFInst_3_n6 ), .B(AddConstOutput[26]), .Z(
        SubCellInst_LFInst_14_LFInst_3_n1 ) );
  AND2 SubCellInst_LFInst_14_LFInst_3_U4  ( .A(AddConstOutput[26]), .B(
        AddConstOutput[25]), .Z(SubCellInst_LFInst_14_LFInst_3_n4 ) );
  ORN2 SubCellInst_LFInst_14_LFInst_3_U3  ( .A(
        SubCellInst_LFInst_14_LFInst_3_n4 ), .B(
        SubCellInst_LFInst_14_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_14_LFInst_3_n3 ) );
  ORN2 SubCellInst_LFInst_14_LFInst_3_U2  ( .A(AddConstOutput[27]), .B(
        SubCellInst_LFInst_14_LFInst_3_n3 ), .Z(
        SubCellInst_LFInst_14_LFInst_3_n2 ) );
  ORN2 SubCellInst_LFInst_14_LFInst_3_U1  ( .A(
        SubCellInst_LFInst_14_LFInst_3_n1 ), .B(
        SubCellInst_LFInst_14_LFInst_3_n2 ), .Z(MCInst1_MC1_v0_3 [0]) );
  BIC2 SubCellInst_LFInst_14_LFInst_2_U11  ( .A(AddConstOutput[25]), .B(
        AddConstOutput[24]), .Z(SubCellInst_LFInst_14_LFInst_2_n8 ) );
  ORN2 SubCellInst_LFInst_14_LFInst_2_U10  ( .A(AddConstOutput[24]), .B(
        AddConstOutput[27]), .Z(SubCellInst_LFInst_14_LFInst_2_n10 ) );
  ORN2 SubCellInst_LFInst_14_LFInst_2_U9  ( .A(AddConstOutput[25]), .B(
        SubCellInst_LFInst_14_LFInst_2_n10 ), .Z(
        SubCellInst_LFInst_14_LFInst_2_n9 ) );
  ORN2 SubCellInst_LFInst_14_LFInst_2_U8  ( .A(
        SubCellInst_LFInst_14_LFInst_2_n8 ), .B(
        SubCellInst_LFInst_14_LFInst_2_n9 ), .Z(
        SubCellInst_LFInst_14_LFInst_2_n7 ) );
  BIC2 SubCellInst_LFInst_14_LFInst_2_U7  ( .A(
        SubCellInst_LFInst_14_LFInst_2_n7 ), .B(AddConstOutput[26]), .Z(
        SubCellInst_LFInst_14_LFInst_2_n1 ) );
  ORN2 SubCellInst_LFInst_14_LFInst_2_U6  ( .A(AddConstOutput[25]), .B(
        AddConstOutput[27]), .Z(SubCellInst_LFInst_14_LFInst_2_n4 ) );
  AND2 SubCellInst_LFInst_14_LFInst_2_U5  ( .A(AddConstOutput[25]), .B(
        AddConstOutput[24]), .Z(SubCellInst_LFInst_14_LFInst_2_n6 ) );
  ORN2 SubCellInst_LFInst_14_LFInst_2_U4  ( .A(AddConstOutput[27]), .B(
        SubCellInst_LFInst_14_LFInst_2_n6 ), .Z(
        SubCellInst_LFInst_14_LFInst_2_n5 ) );
  AND2 SubCellInst_LFInst_14_LFInst_2_U3  ( .A(
        SubCellInst_LFInst_14_LFInst_2_n4 ), .B(
        SubCellInst_LFInst_14_LFInst_2_n5 ), .Z(
        SubCellInst_LFInst_14_LFInst_2_n3 ) );
  ORN2 SubCellInst_LFInst_14_LFInst_2_U2  ( .A(
        SubCellInst_LFInst_14_LFInst_2_n3 ), .B(AddConstOutput[26]), .Z(
        SubCellInst_LFInst_14_LFInst_2_n2 ) );
  ORN2 SubCellInst_LFInst_14_LFInst_2_U1  ( .A(
        SubCellInst_LFInst_14_LFInst_2_n1 ), .B(
        SubCellInst_LFInst_14_LFInst_2_n2 ), .Z(MCInst1_MC1_v0_3 [3]) );
  AND2 SubCellInst_LFInst_14_LFInst_1_U8  ( .A(AddConstOutput[26]), .B(
        AddConstOutput[24]), .Z(SubCellInst_LFInst_14_LFInst_1_n4 ) );
  AND2 SubCellInst_LFInst_14_LFInst_1_U7  ( .A(AddConstOutput[25]), .B(
        AddConstOutput[24]), .Z(SubCellInst_LFInst_14_LFInst_1_n7 ) );
  OR2 SubCellInst_LFInst_14_LFInst_1_U6  ( .A(AddConstOutput[26]), .B(
        SubCellInst_LFInst_14_LFInst_1_n7 ), .Z(
        SubCellInst_LFInst_14_LFInst_1_n6 ) );
  ORN2 SubCellInst_LFInst_14_LFInst_1_U5  ( .A(
        SubCellInst_LFInst_14_LFInst_1_n4 ), .B(
        SubCellInst_LFInst_14_LFInst_1_n6 ), .Z(
        SubCellInst_LFInst_14_LFInst_1_n5 ) );
  AND2 SubCellInst_LFInst_14_LFInst_1_U4  ( .A(AddConstOutput[27]), .B(
        SubCellInst_LFInst_14_LFInst_1_n5 ), .Z(
        SubCellInst_LFInst_14_LFInst_1_n1 ) );
  BIC2 SubCellInst_LFInst_14_LFInst_1_U3  ( .A(AddConstOutput[25]), .B(
        SubCellInst_LFInst_14_LFInst_1_n4 ), .Z(
        SubCellInst_LFInst_14_LFInst_1_n3 ) );
  ORN2 SubCellInst_LFInst_14_LFInst_1_U2  ( .A(AddConstOutput[27]), .B(
        SubCellInst_LFInst_14_LFInst_1_n3 ), .Z(
        SubCellInst_LFInst_14_LFInst_1_n2 ) );
  ORN2 SubCellInst_LFInst_14_LFInst_1_U1  ( .A(
        SubCellInst_LFInst_14_LFInst_1_n1 ), .B(
        SubCellInst_LFInst_14_LFInst_1_n2 ), .Z(MCInst1_MC1_v0_0 [3]) );
  BIC2 SubCellInst_LFInst_14_LFInst_0_U3  ( .A(AddConstOutput[26]), .B(
        AddConstOutput[25]), .Z(SubCellInst_LFInst_14_LFInst_0_n1 ) );
  XOR2 SubCellInst_LFInst_14_LFInst_0_U2  ( .A(AddConstOutput[27]), .B(
        AddConstOutput[24]), .Z(SubCellInst_LFInst_14_LFInst_0_n2 ) );
  XOR2 SubCellInst_LFInst_14_LFInst_0_U1  ( .A(
        SubCellInst_LFInst_14_LFInst_0_n1 ), .B(
        SubCellInst_LFInst_14_LFInst_0_n2 ), .Z(ShiftRowsOutput[56]) );
  OR2 SubCellInst_LFInst_15_LFInst_3_U9  ( .A(AddConstOutput[29]), .B(
        AddConstOutput[28]), .Z(SubCellInst_LFInst_15_LFInst_3_n5 ) );
  AND2 SubCellInst_LFInst_15_LFInst_3_U8  ( .A(AddConstOutput[31]), .B(
        SubCellInst_LFInst_15_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_15_LFInst_3_n7 ) );
  AND2 SubCellInst_LFInst_15_LFInst_3_U7  ( .A(AddConstOutput[28]), .B(
        AddConstOutput[29]), .Z(SubCellInst_LFInst_15_LFInst_3_n8 ) );
  OR2 SubCellInst_LFInst_15_LFInst_3_U6  ( .A(
        SubCellInst_LFInst_15_LFInst_3_n7 ), .B(
        SubCellInst_LFInst_15_LFInst_3_n8 ), .Z(
        SubCellInst_LFInst_15_LFInst_3_n6 ) );
  BIC2 SubCellInst_LFInst_15_LFInst_3_U5  ( .A(
        SubCellInst_LFInst_15_LFInst_3_n6 ), .B(AddConstOutput[30]), .Z(
        SubCellInst_LFInst_15_LFInst_3_n1 ) );
  AND2 SubCellInst_LFInst_15_LFInst_3_U4  ( .A(AddConstOutput[30]), .B(
        AddConstOutput[29]), .Z(SubCellInst_LFInst_15_LFInst_3_n4 ) );
  ORN2 SubCellInst_LFInst_15_LFInst_3_U3  ( .A(
        SubCellInst_LFInst_15_LFInst_3_n4 ), .B(
        SubCellInst_LFInst_15_LFInst_3_n5 ), .Z(
        SubCellInst_LFInst_15_LFInst_3_n3 ) );
  ORN2 SubCellInst_LFInst_15_LFInst_3_U2  ( .A(AddConstOutput[31]), .B(
        SubCellInst_LFInst_15_LFInst_3_n3 ), .Z(
        SubCellInst_LFInst_15_LFInst_3_n2 ) );
  ORN2 SubCellInst_LFInst_15_LFInst_3_U1  ( .A(
        SubCellInst_LFInst_15_LFInst_3_n1 ), .B(
        SubCellInst_LFInst_15_LFInst_3_n2 ), .Z(MCInst1_MC0_v0_3 [0]) );
  BIC2 SubCellInst_LFInst_15_LFInst_2_U11  ( .A(AddConstOutput[29]), .B(
        AddConstOutput[28]), .Z(SubCellInst_LFInst_15_LFInst_2_n8 ) );
  ORN2 SubCellInst_LFInst_15_LFInst_2_U10  ( .A(AddConstOutput[28]), .B(
        AddConstOutput[31]), .Z(SubCellInst_LFInst_15_LFInst_2_n10 ) );
  ORN2 SubCellInst_LFInst_15_LFInst_2_U9  ( .A(AddConstOutput[29]), .B(
        SubCellInst_LFInst_15_LFInst_2_n10 ), .Z(
        SubCellInst_LFInst_15_LFInst_2_n9 ) );
  ORN2 SubCellInst_LFInst_15_LFInst_2_U8  ( .A(
        SubCellInst_LFInst_15_LFInst_2_n8 ), .B(
        SubCellInst_LFInst_15_LFInst_2_n9 ), .Z(
        SubCellInst_LFInst_15_LFInst_2_n7 ) );
  BIC2 SubCellInst_LFInst_15_LFInst_2_U7  ( .A(
        SubCellInst_LFInst_15_LFInst_2_n7 ), .B(AddConstOutput[30]), .Z(
        SubCellInst_LFInst_15_LFInst_2_n1 ) );
  ORN2 SubCellInst_LFInst_15_LFInst_2_U6  ( .A(AddConstOutput[29]), .B(
        AddConstOutput[31]), .Z(SubCellInst_LFInst_15_LFInst_2_n4 ) );
  AND2 SubCellInst_LFInst_15_LFInst_2_U5  ( .A(AddConstOutput[29]), .B(
        AddConstOutput[28]), .Z(SubCellInst_LFInst_15_LFInst_2_n6 ) );
  ORN2 SubCellInst_LFInst_15_LFInst_2_U4  ( .A(AddConstOutput[31]), .B(
        SubCellInst_LFInst_15_LFInst_2_n6 ), .Z(
        SubCellInst_LFInst_15_LFInst_2_n5 ) );
  AND2 SubCellInst_LFInst_15_LFInst_2_U3  ( .A(
        SubCellInst_LFInst_15_LFInst_2_n4 ), .B(
        SubCellInst_LFInst_15_LFInst_2_n5 ), .Z(
        SubCellInst_LFInst_15_LFInst_2_n3 ) );
  ORN2 SubCellInst_LFInst_15_LFInst_2_U2  ( .A(
        SubCellInst_LFInst_15_LFInst_2_n3 ), .B(AddConstOutput[30]), .Z(
        SubCellInst_LFInst_15_LFInst_2_n2 ) );
  ORN2 SubCellInst_LFInst_15_LFInst_2_U1  ( .A(
        SubCellInst_LFInst_15_LFInst_2_n1 ), .B(
        SubCellInst_LFInst_15_LFInst_2_n2 ), .Z(MCInst1_MC0_v0_3 [3]) );
  AND2 SubCellInst_LFInst_15_LFInst_1_U8  ( .A(AddConstOutput[30]), .B(
        AddConstOutput[28]), .Z(SubCellInst_LFInst_15_LFInst_1_n4 ) );
  AND2 SubCellInst_LFInst_15_LFInst_1_U7  ( .A(AddConstOutput[29]), .B(
        AddConstOutput[28]), .Z(SubCellInst_LFInst_15_LFInst_1_n7 ) );
  OR2 SubCellInst_LFInst_15_LFInst_1_U6  ( .A(AddConstOutput[30]), .B(
        SubCellInst_LFInst_15_LFInst_1_n7 ), .Z(
        SubCellInst_LFInst_15_LFInst_1_n6 ) );
  ORN2 SubCellInst_LFInst_15_LFInst_1_U5  ( .A(
        SubCellInst_LFInst_15_LFInst_1_n4 ), .B(
        SubCellInst_LFInst_15_LFInst_1_n6 ), .Z(
        SubCellInst_LFInst_15_LFInst_1_n5 ) );
  AND2 SubCellInst_LFInst_15_LFInst_1_U4  ( .A(AddConstOutput[31]), .B(
        SubCellInst_LFInst_15_LFInst_1_n5 ), .Z(
        SubCellInst_LFInst_15_LFInst_1_n1 ) );
  BIC2 SubCellInst_LFInst_15_LFInst_1_U3  ( .A(AddConstOutput[29]), .B(
        SubCellInst_LFInst_15_LFInst_1_n4 ), .Z(
        SubCellInst_LFInst_15_LFInst_1_n3 ) );
  ORN2 SubCellInst_LFInst_15_LFInst_1_U2  ( .A(AddConstOutput[31]), .B(
        SubCellInst_LFInst_15_LFInst_1_n3 ), .Z(
        SubCellInst_LFInst_15_LFInst_1_n2 ) );
  ORN2 SubCellInst_LFInst_15_LFInst_1_U1  ( .A(
        SubCellInst_LFInst_15_LFInst_1_n1 ), .B(
        SubCellInst_LFInst_15_LFInst_1_n2 ), .Z(MCInst1_MC0_v0_0 [3]) );
  BIC2 SubCellInst_LFInst_15_LFInst_0_U3  ( .A(AddConstOutput[30]), .B(
        AddConstOutput[29]), .Z(SubCellInst_LFInst_15_LFInst_0_n1 ) );
  XOR2 SubCellInst_LFInst_15_LFInst_0_U2  ( .A(AddConstOutput[31]), .B(
        AddConstOutput[28]), .Z(SubCellInst_LFInst_15_LFInst_0_n2 ) );
  XOR2 SubCellInst_LFInst_15_LFInst_0_U1  ( .A(
        SubCellInst_LFInst_15_LFInst_0_n1 ), .B(
        SubCellInst_LFInst_15_LFInst_0_n2 ), .Z(ShiftRowsOutput[60]) );
  XOR2 MCInst1_MC0_v0_2Inst_0_U2  ( .A(MCInst1_MC0_v0_3 [0]), .B(
        MCInst1_MC0_v0_0 [3]), .Z(MCInst1_MC0_v0_2Inst_0_n1 ) );
  XOR2 MCInst1_MC0_v0_2Inst_0_U1  ( .A(ShiftRowsOutput[60]), .B(
        MCInst1_MC0_v0_2Inst_0_n1 ), .Z(MCInst1_MC0_v0_2 [0]) );
  XOR2 MCInst1_MC0_v1_1Inst_0_U1  ( .A(MCInst1_MC0_v1_3 [0]), .B(
        MCInst1_MC0_v1_3 [3]), .Z(MCInst1_MC0_v1_1 [0]) );
  XOR2 MCInst1_MC0_v1_2Inst_0_U2  ( .A(MCInst1_MC0_v1_3 [0]), .B(
        MCInst1_MC0_v1_3 [3]), .Z(MCInst1_MC0_v1_2Inst_0_n1 ) );
  XOR2 MCInst1_MC0_v1_2Inst_0_U1  ( .A(MCInst1_MC0_v1_3 [2]), .B(
        MCInst1_MC0_v1_2Inst_0_n1 ), .Z(MCInst1_MC0_v1_2 [0]) );
  XOR2 MCInst1_MC0_v2_1Inst_0_U1  ( .A(MCInst1_MC0_v2_0 [3]), .B(
        MCInst1_MC0_v2_3 [1]), .Z(MCInst1_MC0_v2_1 [0]) );
  XOR2 MCInst1_MC0_v2_2Inst_0_U1  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v2_0 [2]), .Z(MCInst1_MC0_v2_2 [0]) );
  XOR2 MCInst1_MC0_v2_3Inst_0_U3  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v2_0 [3]), .Z(MCInst1_MC0_v2_3Inst_0_n1 ) );
  XOR2 MCInst1_MC0_v2_3Inst_0_U2  ( .A(MCInst1_MC0_v2_0 [2]), .B(
        MCInst1_MC0_v2_3 [1]), .Z(MCInst1_MC0_v2_3Inst_0_n2 ) );
  XOR2 MCInst1_MC0_v2_3Inst_0_U1  ( .A(MCInst1_MC0_v2_3Inst_0_n1 ), .B(
        MCInst1_MC0_v2_3Inst_0_n2 ), .Z(MCInst1_MC0_v2_3 [0]) );
  XOR2 MCInst1_MC0_v3_1Inst_0_U1  ( .A(MCInst1_MC0_v3_2 [2]), .B(
        MCInst1_MC0_v3_0 [3]), .Z(MCInst1_MC0_v3_1 [0]) );
  XOR2 MCInst1_MC0_v3_2Inst_0_U1  ( .A(MCInst1_MC0_v3_0 [2]), .B(
        MCInst1_MC0_v3_2 [3]), .Z(MCInst1_MC0_v3_2 [0]) );
  XOR2 MCInst1_MC0_v3_3Inst_0_U2  ( .A(MCInst1_MC0_v3_2 [2]), .B(
        MCInst1_MC0_v3_0 [2]), .Z(MCInst1_MC0_v3_3Inst_0_n1 ) );
  XOR2 MCInst1_MC0_v3_3Inst_0_U1  ( .A(MCInst1_MC0_v3_2 [3]), .B(
        MCInst1_MC0_v3_3Inst_0_n1 ), .Z(MCInst1_MC0_v3_3 [0]) );
  XOR2 MCInst1_MC0_v0_0Inst_1_U1  ( .A(MCInst1_MC0_v0_3 [0]), .B(
        MCInst1_MC0_v0_3 [3]), .Z(MCInst1_MC0_v0_0 [1]) );
  XOR2 MCInst1_MC0_v0_1Inst_1_U1  ( .A(MCInst1_MC0_v0_3 [3]), .B(
        MCInst1_MC0_v0_0 [3]), .Z(MCInst1_MC0_v0_1 [1]) );
  XOR2 MCInst1_MC0_v0_2Inst_1_U2  ( .A(MCInst1_MC0_v0_3 [0]), .B(
        MCInst1_MC0_v0_3 [3]), .Z(MCInst1_MC0_v0_2Inst_1_n1 ) );
  XOR2 MCInst1_MC0_v0_2Inst_1_U1  ( .A(ShiftRowsOutput[60]), .B(
        MCInst1_MC0_v0_2Inst_1_n1 ), .Z(MCInst1_MC0_v0_2 [1]) );
  XOR2 MCInst1_MC0_v0_3Inst_1_U1  ( .A(MCInst1_MC0_v0_3 [0]), .B(
        ShiftRowsOutput[60]), .Z(MCInst1_MC0_v0_3 [1]) );
  XOR2 MCInst1_MC0_v1_1Inst_1_U1  ( .A(MCInst1_MC0_v1_3 [3]), .B(
        ShiftRowsOutput[44]), .Z(MCInst1_MC0_v1_1 [1]) );
  XOR2 MCInst1_MC0_v1_2Inst_1_U1  ( .A(MCInst1_MC0_v1_3 [2]), .B(
        ShiftRowsOutput[44]), .Z(MCInst1_MC0_v1_2 [1]) );
  XOR2 MCInst1_MC0_v1_3Inst_1_U1  ( .A(MCInst1_MC0_v1_3 [0]), .B(
        ShiftRowsOutput[44]), .Z(MCInst1_MC0_v1_3 [1]) );
  XOR2 MCInst1_MC0_v2_0Inst_1_U1  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v2_3 [1]), .Z(MCInst1_MC0_v2_0 [1]) );
  XOR2 MCInst1_MC0_v2_1Inst_1_U2  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v2_0 [3]), .Z(MCInst1_MC0_v2_1Inst_1_n1 ) );
  XOR2 MCInst1_MC0_v2_1Inst_1_U1  ( .A(MCInst1_MC0_v2_0 [2]), .B(
        MCInst1_MC0_v2_1Inst_1_n1 ), .Z(MCInst1_MC0_v2_1 [1]) );
  XOR2 MCInst1_MC0_v2_2Inst_1_U3  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v2_0 [3]), .Z(MCInst1_MC0_v2_2Inst_1_n1 ) );
  XOR2 MCInst1_MC0_v2_2Inst_1_U2  ( .A(MCInst1_MC0_v2_0 [2]), .B(
        MCInst1_MC0_v2_3 [1]), .Z(MCInst1_MC0_v2_2Inst_1_n2 ) );
  XOR2 MCInst1_MC0_v2_2Inst_1_U1  ( .A(MCInst1_MC0_v2_2Inst_1_n1 ), .B(
        MCInst1_MC0_v2_2Inst_1_n2 ), .Z(MCInst1_MC0_v2_2 [1]) );
  XOR2 MCInst1_MC0_v3_0Inst_1_U1  ( .A(MCInst1_MC0_v3_2 [2]), .B(
        MCInst1_MC0_v3_2 [3]), .Z(MCInst1_MC0_v3_0 [1]) );
  XOR2 MCInst1_MC0_v3_1Inst_1_U1  ( .A(MCInst1_MC0_v3_0 [3]), .B(
        MCInst1_MC0_v3_2 [3]), .Z(MCInst1_MC0_v3_1 [1]) );
  XOR2 MCInst1_MC0_v3_3Inst_1_U2  ( .A(MCInst1_MC0_v3_2 [2]), .B(
        MCInst1_MC0_v3_0 [3]), .Z(MCInst1_MC0_v3_3Inst_1_n1 ) );
  XOR2 MCInst1_MC0_v3_3Inst_1_U1  ( .A(MCInst1_MC0_v3_2 [3]), .B(
        MCInst1_MC0_v3_3Inst_1_n1 ), .Z(MCInst1_MC0_v3_3 [1]) );
  XOR2 MCInst1_MC0_v0_0Inst_2_U1  ( .A(MCInst1_MC0_v0_3 [0]), .B(
        ShiftRowsOutput[60]), .Z(MCInst1_MC0_v0_0 [2]) );
  XOR2 MCInst1_MC0_v0_1Inst_2_U1  ( .A(MCInst1_MC0_v0_3 [0]), .B(
        MCInst1_MC0_v0_3 [3]), .Z(MCInst1_MC0_v0_1 [2]) );
  XOR2 MCInst1_MC0_v0_2Inst_2_U1  ( .A(MCInst1_MC0_v0_3 [0]), .B(
        MCInst1_MC0_v0_0 [3]), .Z(MCInst1_MC0_v0_2 [2]) );
  XOR2 MCInst1_MC0_v1_1Inst_2_U2  ( .A(MCInst1_MC0_v1_3 [0]), .B(
        MCInst1_MC0_v1_3 [2]), .Z(MCInst1_MC0_v1_1Inst_2_n1 ) );
  XOR2 MCInst1_MC0_v1_1Inst_2_U1  ( .A(ShiftRowsOutput[44]), .B(
        MCInst1_MC0_v1_1Inst_2_n1 ), .Z(MCInst1_MC0_v1_1 [2]) );
  XOR2 MCInst1_MC0_v1_2Inst_2_U2  ( .A(MCInst1_MC0_v1_3 [3]), .B(
        MCInst1_MC0_v1_3 [2]), .Z(MCInst1_MC0_v1_2Inst_2_n1 ) );
  XOR2 MCInst1_MC0_v1_2Inst_2_U1  ( .A(ShiftRowsOutput[44]), .B(
        MCInst1_MC0_v1_2Inst_2_n1 ), .Z(MCInst1_MC0_v1_2 [2]) );
  XOR2 MCInst1_MC0_v2_1Inst_2_U2  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v2_0 [3]), .Z(MCInst1_MC0_v2_1Inst_2_n1 ) );
  XOR2 MCInst1_MC0_v2_1Inst_2_U1  ( .A(MCInst1_MC0_v2_3 [1]), .B(
        MCInst1_MC0_v2_1Inst_2_n1 ), .Z(MCInst1_MC0_v2_1 [2]) );
  XOR2 MCInst1_MC0_v2_2Inst_2_U2  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v2_0 [3]), .Z(MCInst1_MC0_v2_2Inst_2_n1 ) );
  XOR2 MCInst1_MC0_v2_2Inst_2_U1  ( .A(MCInst1_MC0_v2_0 [2]), .B(
        MCInst1_MC0_v2_2Inst_2_n1 ), .Z(MCInst1_MC0_v2_2 [2]) );
  XOR2 MCInst1_MC0_v2_3Inst_2_U1  ( .A(MCInst1_MC0_v2_0 [2]), .B(
        MCInst1_MC0_v2_3 [1]), .Z(MCInst1_MC0_v2_3 [2]) );
  XOR2 MCInst1_MC0_v3_1Inst_2_U2  ( .A(MCInst1_MC0_v3_2 [2]), .B(
        MCInst1_MC0_v3_0 [2]), .Z(MCInst1_MC0_v3_1Inst_2_n1 ) );
  XOR2 MCInst1_MC0_v3_1Inst_2_U1  ( .A(MCInst1_MC0_v3_2 [3]), .B(
        MCInst1_MC0_v3_1Inst_2_n1 ), .Z(MCInst1_MC0_v3_1 [2]) );
  XOR2 MCInst1_MC0_v3_3Inst_2_U1  ( .A(MCInst1_MC0_v3_2 [2]), .B(
        MCInst1_MC0_v3_0 [2]), .Z(MCInst1_MC0_v3_3 [2]) );
  XOR2 MCInst1_MC0_v0_1Inst_3_U1  ( .A(MCInst1_MC0_v0_3 [0]), .B(
        ShiftRowsOutput[60]), .Z(MCInst1_MC0_v0_1 [3]) );
  XOR2 MCInst1_MC0_v0_2Inst_3_U1  ( .A(MCInst1_MC0_v0_3 [3]), .B(
        ShiftRowsOutput[60]), .Z(MCInst1_MC0_v0_2 [3]) );
  XOR2 MCInst1_MC0_v1_1Inst_3_U1  ( .A(MCInst1_MC0_v1_3 [3]), .B(
        MCInst1_MC0_v1_3 [2]), .Z(MCInst1_MC0_v1_1 [3]) );
  XOR2 MCInst1_MC0_v1_2Inst_3_U3  ( .A(MCInst1_MC0_v1_3 [0]), .B(
        MCInst1_MC0_v1_3 [3]), .Z(MCInst1_MC0_v1_2Inst_3_n1 ) );
  XOR2 MCInst1_MC0_v1_2Inst_3_U2  ( .A(MCInst1_MC0_v1_3 [2]), .B(
        ShiftRowsOutput[44]), .Z(MCInst1_MC0_v1_2Inst_3_n2 ) );
  XOR2 MCInst1_MC0_v1_2Inst_3_U1  ( .A(MCInst1_MC0_v1_2Inst_3_n1 ), .B(
        MCInst1_MC0_v1_2Inst_3_n2 ), .Z(MCInst1_MC0_v1_2 [3]) );
  XOR2 MCInst1_MC0_v2_1Inst_3_U1  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v2_0 [2]), .Z(MCInst1_MC0_v2_1 [3]) );
  XOR2 MCInst1_MC0_v2_2Inst_3_U2  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v2_0 [3]), .Z(MCInst1_MC0_v2_2Inst_3_n1 ) );
  XOR2 MCInst1_MC0_v2_2Inst_3_U1  ( .A(MCInst1_MC0_v2_3 [1]), .B(
        MCInst1_MC0_v2_2Inst_3_n1 ), .Z(MCInst1_MC0_v2_2 [3]) );
  XOR2 MCInst1_MC0_v2_3Inst_3_U2  ( .A(MCInst1_MC0_v2_0 [3]), .B(
        MCInst1_MC0_v2_0 [2]), .Z(MCInst1_MC0_v2_3Inst_3_n1 ) );
  XOR2 MCInst1_MC0_v2_3Inst_3_U1  ( .A(MCInst1_MC0_v2_3 [1]), .B(
        MCInst1_MC0_v2_3Inst_3_n1 ), .Z(MCInst1_MC0_v2_3 [3]) );
  XOR2 MCInst1_MC0_v3_1Inst_3_U1  ( .A(MCInst1_MC0_v3_0 [3]), .B(
        MCInst1_MC0_v3_0 [2]), .Z(MCInst1_MC0_v3_1 [3]) );
  XOR2 MCInst1_MC0_v3_3Inst_3_U1  ( .A(MCInst1_MC0_v3_0 [3]), .B(
        MCInst1_MC0_v3_2 [3]), .Z(MCInst1_MC0_v3_3 [3]) );
  XOR2 MCInst1_MC0_r0Inst_XORInst_0_0_U4  ( .A(
        MCInst1_MC0_r0Inst_XORInst_0_0_n2 ), .B(
        MCInst1_MC0_r0Inst_XORInst_0_0_n1 ), .Z(Feedback[60]) );
  XOR2 MCInst1_MC0_r0Inst_XORInst_0_0_U3  ( .A(1'b0), .B(
        MCInst1_MC0_r0Inst_XORInst_0_0_n3 ), .Z(
        MCInst1_MC0_r0Inst_XORInst_0_0_n1 ) );
  XOR2 MCInst1_MC0_r0Inst_XORInst_0_0_U2  ( .A(MCInst1_MC0_v2_0 [0]), .B(
        MCInst1_MC0_v3_2 [2]), .Z(MCInst1_MC0_r0Inst_XORInst_0_0_n2 ) );
  XOR2 MCInst1_MC0_r0Inst_XORInst_0_0_U1  ( .A(MCInst1_MC0_v0_3 [3]), .B(
        ShiftRowsOutput[44]), .Z(MCInst1_MC0_r0Inst_XORInst_0_0_n3 ) );
  XOR2 MCInst1_MC0_r0Inst_XORInst_0_1_U4  ( .A(
        MCInst1_MC0_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC0_r0Inst_XORInst_0_1_n6 ), .Z(Feedback[61]) );
  XOR2 MCInst1_MC0_r0Inst_XORInst_0_1_U3  ( .A(1'b0), .B(
        MCInst1_MC0_r0Inst_XORInst_0_1_n4 ), .Z(
        MCInst1_MC0_r0Inst_XORInst_0_1_n6 ) );
  XOR2 MCInst1_MC0_r0Inst_XORInst_0_1_U2  ( .A(MCInst1_MC0_v2_0 [1]), .B(
        MCInst1_MC0_v3_0 [1]), .Z(MCInst1_MC0_r0Inst_XORInst_0_1_n5 ) );
  XOR2 MCInst1_MC0_r0Inst_XORInst_0_1_U1  ( .A(MCInst1_MC0_v0_0 [1]), .B(
        MCInst1_MC0_v1_3 [2]), .Z(MCInst1_MC0_r0Inst_XORInst_0_1_n4 ) );
  XOR2 MCInst1_MC0_r0Inst_XORInst_0_2_U4  ( .A(
        MCInst1_MC0_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC0_r0Inst_XORInst_0_2_n6 ), .Z(Feedback[62]) );
  XOR2 MCInst1_MC0_r0Inst_XORInst_0_2_U3  ( .A(1'b0), .B(
        MCInst1_MC0_r0Inst_XORInst_0_2_n4 ), .Z(
        MCInst1_MC0_r0Inst_XORInst_0_2_n6 ) );
  XOR2 MCInst1_MC0_r0Inst_XORInst_0_2_U2  ( .A(MCInst1_MC0_v2_0 [2]), .B(
        MCInst1_MC0_v3_0 [2]), .Z(MCInst1_MC0_r0Inst_XORInst_0_2_n5 ) );
  XOR2 MCInst1_MC0_r0Inst_XORInst_0_2_U1  ( .A(MCInst1_MC0_v0_0 [2]), .B(
        MCInst1_MC0_v1_3 [3]), .Z(MCInst1_MC0_r0Inst_XORInst_0_2_n4 ) );
  XOR2 MCInst1_MC0_r0Inst_XORInst_0_3_U4  ( .A(
        MCInst1_MC0_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC0_r0Inst_XORInst_0_3_n6 ), .Z(Feedback[63]) );
  XOR2 MCInst1_MC0_r0Inst_XORInst_0_3_U3  ( .A(1'b0), .B(
        MCInst1_MC0_r0Inst_XORInst_0_3_n4 ), .Z(
        MCInst1_MC0_r0Inst_XORInst_0_3_n6 ) );
  XOR2 MCInst1_MC0_r0Inst_XORInst_0_3_U2  ( .A(MCInst1_MC0_v2_0 [3]), .B(
        MCInst1_MC0_v3_0 [3]), .Z(MCInst1_MC0_r0Inst_XORInst_0_3_n5 ) );
  XOR2 MCInst1_MC0_r0Inst_XORInst_0_3_U1  ( .A(MCInst1_MC0_v0_0 [3]), .B(
        MCInst1_MC0_v1_3 [0]), .Z(MCInst1_MC0_r0Inst_XORInst_0_3_n4 ) );
  XOR2 MCInst1_MC0_r1Inst_XORInst_0_0_U4  ( .A(
        MCInst1_MC0_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC0_r1Inst_XORInst_0_0_n6 ), .Z(Feedback[44]) );
  XOR2 MCInst1_MC0_r1Inst_XORInst_0_0_U3  ( .A(1'b0), .B(
        MCInst1_MC0_r1Inst_XORInst_0_0_n4 ), .Z(
        MCInst1_MC0_r1Inst_XORInst_0_0_n6 ) );
  XOR2 MCInst1_MC0_r1Inst_XORInst_0_0_U2  ( .A(MCInst1_MC0_v2_1 [0]), .B(
        MCInst1_MC0_v3_1 [0]), .Z(MCInst1_MC0_r1Inst_XORInst_0_0_n5 ) );
  XOR2 MCInst1_MC0_r1Inst_XORInst_0_0_U1  ( .A(MCInst1_MC0_v0_0 [3]), .B(
        MCInst1_MC0_v1_1 [0]), .Z(MCInst1_MC0_r1Inst_XORInst_0_0_n4 ) );
  XOR2 MCInst1_MC0_r1Inst_XORInst_0_1_U4  ( .A(
        MCInst1_MC0_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC0_r1Inst_XORInst_0_1_n6 ), .Z(Feedback[45]) );
  XOR2 MCInst1_MC0_r1Inst_XORInst_0_1_U3  ( .A(1'b0), .B(
        MCInst1_MC0_r1Inst_XORInst_0_1_n4 ), .Z(
        MCInst1_MC0_r1Inst_XORInst_0_1_n6 ) );
  XOR2 MCInst1_MC0_r1Inst_XORInst_0_1_U2  ( .A(MCInst1_MC0_v2_1 [1]), .B(
        MCInst1_MC0_v3_1 [1]), .Z(MCInst1_MC0_r1Inst_XORInst_0_1_n5 ) );
  XOR2 MCInst1_MC0_r1Inst_XORInst_0_1_U1  ( .A(MCInst1_MC0_v0_1 [1]), .B(
        MCInst1_MC0_v1_1 [1]), .Z(MCInst1_MC0_r1Inst_XORInst_0_1_n4 ) );
  XOR2 MCInst1_MC0_r1Inst_XORInst_0_2_U4  ( .A(
        MCInst1_MC0_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC0_r1Inst_XORInst_0_2_n6 ), .Z(Feedback[46]) );
  XOR2 MCInst1_MC0_r1Inst_XORInst_0_2_U3  ( .A(1'b0), .B(
        MCInst1_MC0_r1Inst_XORInst_0_2_n4 ), .Z(
        MCInst1_MC0_r1Inst_XORInst_0_2_n6 ) );
  XOR2 MCInst1_MC0_r1Inst_XORInst_0_2_U2  ( .A(MCInst1_MC0_v2_1 [2]), .B(
        MCInst1_MC0_v3_1 [2]), .Z(MCInst1_MC0_r1Inst_XORInst_0_2_n5 ) );
  XOR2 MCInst1_MC0_r1Inst_XORInst_0_2_U1  ( .A(MCInst1_MC0_v0_1 [2]), .B(
        MCInst1_MC0_v1_1 [2]), .Z(MCInst1_MC0_r1Inst_XORInst_0_2_n4 ) );
  XOR2 MCInst1_MC0_r1Inst_XORInst_0_3_U4  ( .A(
        MCInst1_MC0_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC0_r1Inst_XORInst_0_3_n6 ), .Z(Feedback[47]) );
  XOR2 MCInst1_MC0_r1Inst_XORInst_0_3_U3  ( .A(1'b0), .B(
        MCInst1_MC0_r1Inst_XORInst_0_3_n4 ), .Z(
        MCInst1_MC0_r1Inst_XORInst_0_3_n6 ) );
  XOR2 MCInst1_MC0_r1Inst_XORInst_0_3_U2  ( .A(MCInst1_MC0_v2_1 [3]), .B(
        MCInst1_MC0_v3_1 [3]), .Z(MCInst1_MC0_r1Inst_XORInst_0_3_n5 ) );
  XOR2 MCInst1_MC0_r1Inst_XORInst_0_3_U1  ( .A(MCInst1_MC0_v0_1 [3]), .B(
        MCInst1_MC0_v1_1 [3]), .Z(MCInst1_MC0_r1Inst_XORInst_0_3_n4 ) );
  XOR2 MCInst1_MC0_r2Inst_XORInst_0_0_U4  ( .A(
        MCInst1_MC0_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC0_r2Inst_XORInst_0_0_n6 ), .Z(Feedback[28]) );
  XOR2 MCInst1_MC0_r2Inst_XORInst_0_0_U3  ( .A(1'b0), .B(
        MCInst1_MC0_r2Inst_XORInst_0_0_n4 ), .Z(
        MCInst1_MC0_r2Inst_XORInst_0_0_n6 ) );
  XOR2 MCInst1_MC0_r2Inst_XORInst_0_0_U2  ( .A(MCInst1_MC0_v2_2 [0]), .B(
        MCInst1_MC0_v3_2 [0]), .Z(MCInst1_MC0_r2Inst_XORInst_0_0_n5 ) );
  XOR2 MCInst1_MC0_r2Inst_XORInst_0_0_U1  ( .A(MCInst1_MC0_v0_2 [0]), .B(
        MCInst1_MC0_v1_2 [0]), .Z(MCInst1_MC0_r2Inst_XORInst_0_0_n4 ) );
  XOR2 MCInst1_MC0_r2Inst_XORInst_0_1_U4  ( .A(
        MCInst1_MC0_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC0_r2Inst_XORInst_0_1_n6 ), .Z(Feedback[29]) );
  XOR2 MCInst1_MC0_r2Inst_XORInst_0_1_U3  ( .A(1'b0), .B(
        MCInst1_MC0_r2Inst_XORInst_0_1_n4 ), .Z(
        MCInst1_MC0_r2Inst_XORInst_0_1_n6 ) );
  XOR2 MCInst1_MC0_r2Inst_XORInst_0_1_U2  ( .A(MCInst1_MC0_v2_2 [1]), .B(
        MCInst1_MC0_v3_0 [3]), .Z(MCInst1_MC0_r2Inst_XORInst_0_1_n5 ) );
  XOR2 MCInst1_MC0_r2Inst_XORInst_0_1_U1  ( .A(MCInst1_MC0_v0_2 [1]), .B(
        MCInst1_MC0_v1_2 [1]), .Z(MCInst1_MC0_r2Inst_XORInst_0_1_n4 ) );
  XOR2 MCInst1_MC0_r2Inst_XORInst_0_2_U4  ( .A(
        MCInst1_MC0_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC0_r2Inst_XORInst_0_2_n6 ), .Z(Feedback[30]) );
  XOR2 MCInst1_MC0_r2Inst_XORInst_0_2_U3  ( .A(1'b0), .B(
        MCInst1_MC0_r2Inst_XORInst_0_2_n4 ), .Z(
        MCInst1_MC0_r2Inst_XORInst_0_2_n6 ) );
  XOR2 MCInst1_MC0_r2Inst_XORInst_0_2_U2  ( .A(MCInst1_MC0_v2_2 [2]), .B(
        MCInst1_MC0_v3_2 [2]), .Z(MCInst1_MC0_r2Inst_XORInst_0_2_n5 ) );
  XOR2 MCInst1_MC0_r2Inst_XORInst_0_2_U1  ( .A(MCInst1_MC0_v0_2 [2]), .B(
        MCInst1_MC0_v1_2 [2]), .Z(MCInst1_MC0_r2Inst_XORInst_0_2_n4 ) );
  XOR2 MCInst1_MC0_r2Inst_XORInst_0_3_U4  ( .A(
        MCInst1_MC0_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC0_r2Inst_XORInst_0_3_n6 ), .Z(Feedback[31]) );
  XOR2 MCInst1_MC0_r2Inst_XORInst_0_3_U3  ( .A(1'b0), .B(
        MCInst1_MC0_r2Inst_XORInst_0_3_n4 ), .Z(
        MCInst1_MC0_r2Inst_XORInst_0_3_n6 ) );
  XOR2 MCInst1_MC0_r2Inst_XORInst_0_3_U2  ( .A(MCInst1_MC0_v2_2 [3]), .B(
        MCInst1_MC0_v3_2 [3]), .Z(MCInst1_MC0_r2Inst_XORInst_0_3_n5 ) );
  XOR2 MCInst1_MC0_r2Inst_XORInst_0_3_U1  ( .A(MCInst1_MC0_v0_2 [3]), .B(
        MCInst1_MC0_v1_2 [3]), .Z(MCInst1_MC0_r2Inst_XORInst_0_3_n4 ) );
  XOR2 MCInst1_MC0_r3Inst_XORInst_0_0_U4  ( .A(
        MCInst1_MC0_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC0_r3Inst_XORInst_0_0_n6 ), .Z(Feedback[12]) );
  XOR2 MCInst1_MC0_r3Inst_XORInst_0_0_U3  ( .A(1'b0), .B(
        MCInst1_MC0_r3Inst_XORInst_0_0_n4 ), .Z(
        MCInst1_MC0_r3Inst_XORInst_0_0_n6 ) );
  XOR2 MCInst1_MC0_r3Inst_XORInst_0_0_U2  ( .A(MCInst1_MC0_v2_3 [0]), .B(
        MCInst1_MC0_v3_3 [0]), .Z(MCInst1_MC0_r3Inst_XORInst_0_0_n5 ) );
  XOR2 MCInst1_MC0_r3Inst_XORInst_0_0_U1  ( .A(MCInst1_MC0_v0_3 [0]), .B(
        MCInst1_MC0_v1_3 [0]), .Z(MCInst1_MC0_r3Inst_XORInst_0_0_n4 ) );
  XOR2 MCInst1_MC0_r3Inst_XORInst_0_1_U4  ( .A(
        MCInst1_MC0_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC0_r3Inst_XORInst_0_1_n6 ), .Z(Feedback[13]) );
  XOR2 MCInst1_MC0_r3Inst_XORInst_0_1_U3  ( .A(1'b0), .B(
        MCInst1_MC0_r3Inst_XORInst_0_1_n4 ), .Z(
        MCInst1_MC0_r3Inst_XORInst_0_1_n6 ) );
  XOR2 MCInst1_MC0_r3Inst_XORInst_0_1_U2  ( .A(MCInst1_MC0_v2_3 [1]), .B(
        MCInst1_MC0_v3_3 [1]), .Z(MCInst1_MC0_r3Inst_XORInst_0_1_n5 ) );
  XOR2 MCInst1_MC0_r3Inst_XORInst_0_1_U1  ( .A(MCInst1_MC0_v0_3 [1]), .B(
        MCInst1_MC0_v1_3 [1]), .Z(MCInst1_MC0_r3Inst_XORInst_0_1_n4 ) );
  XOR2 MCInst1_MC0_r3Inst_XORInst_0_2_U4  ( .A(
        MCInst1_MC0_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC0_r3Inst_XORInst_0_2_n6 ), .Z(Feedback[14]) );
  XOR2 MCInst1_MC0_r3Inst_XORInst_0_2_U3  ( .A(1'b0), .B(
        MCInst1_MC0_r3Inst_XORInst_0_2_n4 ), .Z(
        MCInst1_MC0_r3Inst_XORInst_0_2_n6 ) );
  XOR2 MCInst1_MC0_r3Inst_XORInst_0_2_U2  ( .A(MCInst1_MC0_v2_3 [2]), .B(
        MCInst1_MC0_v3_3 [2]), .Z(MCInst1_MC0_r3Inst_XORInst_0_2_n5 ) );
  XOR2 MCInst1_MC0_r3Inst_XORInst_0_2_U1  ( .A(MCInst1_MC0_v0_0 [3]), .B(
        MCInst1_MC0_v1_3 [2]), .Z(MCInst1_MC0_r3Inst_XORInst_0_2_n4 ) );
  XOR2 MCInst1_MC0_r3Inst_XORInst_0_3_U4  ( .A(
        MCInst1_MC0_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC0_r3Inst_XORInst_0_3_n6 ), .Z(Feedback[15]) );
  XOR2 MCInst1_MC0_r3Inst_XORInst_0_3_U3  ( .A(1'b0), .B(
        MCInst1_MC0_r3Inst_XORInst_0_3_n4 ), .Z(
        MCInst1_MC0_r3Inst_XORInst_0_3_n6 ) );
  XOR2 MCInst1_MC0_r3Inst_XORInst_0_3_U2  ( .A(MCInst1_MC0_v2_3 [3]), .B(
        MCInst1_MC0_v3_3 [3]), .Z(MCInst1_MC0_r3Inst_XORInst_0_3_n5 ) );
  XOR2 MCInst1_MC0_r3Inst_XORInst_0_3_U1  ( .A(MCInst1_MC0_v0_3 [3]), .B(
        MCInst1_MC0_v1_3 [3]), .Z(MCInst1_MC0_r3Inst_XORInst_0_3_n4 ) );
  XOR2 MCInst1_MC1_v0_2Inst_0_U2  ( .A(MCInst1_MC1_v0_3 [0]), .B(
        MCInst1_MC1_v0_0 [3]), .Z(MCInst1_MC1_v0_2Inst_0_n1 ) );
  XOR2 MCInst1_MC1_v0_2Inst_0_U1  ( .A(ShiftRowsOutput[56]), .B(
        MCInst1_MC1_v0_2Inst_0_n1 ), .Z(MCInst1_MC1_v0_2 [0]) );
  XOR2 MCInst1_MC1_v1_1Inst_0_U1  ( .A(MCInst1_MC1_v1_3 [0]), .B(
        MCInst1_MC1_v1_3 [3]), .Z(MCInst1_MC1_v1_1 [0]) );
  XOR2 MCInst1_MC1_v1_2Inst_0_U2  ( .A(MCInst1_MC1_v1_3 [0]), .B(
        MCInst1_MC1_v1_3 [3]), .Z(MCInst1_MC1_v1_2Inst_0_n1 ) );
  XOR2 MCInst1_MC1_v1_2Inst_0_U1  ( .A(MCInst1_MC1_v1_3 [2]), .B(
        MCInst1_MC1_v1_2Inst_0_n1 ), .Z(MCInst1_MC1_v1_2 [0]) );
  XOR2 MCInst1_MC1_v2_1Inst_0_U1  ( .A(MCInst1_MC1_v2_0 [3]), .B(
        MCInst1_MC1_v2_3 [1]), .Z(MCInst1_MC1_v2_1 [0]) );
  XOR2 MCInst1_MC1_v2_2Inst_0_U1  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v2_0 [2]), .Z(MCInst1_MC1_v2_2 [0]) );
  XOR2 MCInst1_MC1_v2_3Inst_0_U3  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v2_0 [3]), .Z(MCInst1_MC1_v2_3Inst_0_n1 ) );
  XOR2 MCInst1_MC1_v2_3Inst_0_U2  ( .A(MCInst1_MC1_v2_0 [2]), .B(
        MCInst1_MC1_v2_3 [1]), .Z(MCInst1_MC1_v2_3Inst_0_n2 ) );
  XOR2 MCInst1_MC1_v2_3Inst_0_U1  ( .A(MCInst1_MC1_v2_3Inst_0_n1 ), .B(
        MCInst1_MC1_v2_3Inst_0_n2 ), .Z(MCInst1_MC1_v2_3 [0]) );
  XOR2 MCInst1_MC1_v3_1Inst_0_U1  ( .A(MCInst1_MC1_v3_2 [2]), .B(
        MCInst1_MC1_v3_0 [3]), .Z(MCInst1_MC1_v3_1 [0]) );
  XOR2 MCInst1_MC1_v3_2Inst_0_U1  ( .A(MCInst1_MC1_v3_0 [2]), .B(
        MCInst1_MC1_v3_2 [3]), .Z(MCInst1_MC1_v3_2 [0]) );
  XOR2 MCInst1_MC1_v3_3Inst_0_U2  ( .A(MCInst1_MC1_v3_2 [2]), .B(
        MCInst1_MC1_v3_0 [2]), .Z(MCInst1_MC1_v3_3Inst_0_n1 ) );
  XOR2 MCInst1_MC1_v3_3Inst_0_U1  ( .A(MCInst1_MC1_v3_2 [3]), .B(
        MCInst1_MC1_v3_3Inst_0_n1 ), .Z(MCInst1_MC1_v3_3 [0]) );
  XOR2 MCInst1_MC1_v0_0Inst_1_U1  ( .A(MCInst1_MC1_v0_3 [0]), .B(
        MCInst1_MC1_v0_3 [3]), .Z(MCInst1_MC1_v0_0 [1]) );
  XOR2 MCInst1_MC1_v0_1Inst_1_U1  ( .A(MCInst1_MC1_v0_3 [3]), .B(
        MCInst1_MC1_v0_0 [3]), .Z(MCInst1_MC1_v0_1 [1]) );
  XOR2 MCInst1_MC1_v0_2Inst_1_U2  ( .A(MCInst1_MC1_v0_3 [0]), .B(
        MCInst1_MC1_v0_3 [3]), .Z(MCInst1_MC1_v0_2Inst_1_n1 ) );
  XOR2 MCInst1_MC1_v0_2Inst_1_U1  ( .A(ShiftRowsOutput[56]), .B(
        MCInst1_MC1_v0_2Inst_1_n1 ), .Z(MCInst1_MC1_v0_2 [1]) );
  XOR2 MCInst1_MC1_v0_3Inst_1_U1  ( .A(MCInst1_MC1_v0_3 [0]), .B(
        ShiftRowsOutput[56]), .Z(MCInst1_MC1_v0_3 [1]) );
  XOR2 MCInst1_MC1_v1_1Inst_1_U1  ( .A(MCInst1_MC1_v1_3 [3]), .B(
        ShiftRowsOutput[40]), .Z(MCInst1_MC1_v1_1 [1]) );
  XOR2 MCInst1_MC1_v1_2Inst_1_U1  ( .A(MCInst1_MC1_v1_3 [2]), .B(
        ShiftRowsOutput[40]), .Z(MCInst1_MC1_v1_2 [1]) );
  XOR2 MCInst1_MC1_v1_3Inst_1_U1  ( .A(MCInst1_MC1_v1_3 [0]), .B(
        ShiftRowsOutput[40]), .Z(MCInst1_MC1_v1_3 [1]) );
  XOR2 MCInst1_MC1_v2_0Inst_1_U1  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v2_3 [1]), .Z(MCInst1_MC1_v2_0 [1]) );
  XOR2 MCInst1_MC1_v2_1Inst_1_U2  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v2_0 [3]), .Z(MCInst1_MC1_v2_1Inst_1_n1 ) );
  XOR2 MCInst1_MC1_v2_1Inst_1_U1  ( .A(MCInst1_MC1_v2_0 [2]), .B(
        MCInst1_MC1_v2_1Inst_1_n1 ), .Z(MCInst1_MC1_v2_1 [1]) );
  XOR2 MCInst1_MC1_v2_2Inst_1_U3  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v2_0 [3]), .Z(MCInst1_MC1_v2_2Inst_1_n1 ) );
  XOR2 MCInst1_MC1_v2_2Inst_1_U2  ( .A(MCInst1_MC1_v2_0 [2]), .B(
        MCInst1_MC1_v2_3 [1]), .Z(MCInst1_MC1_v2_2Inst_1_n2 ) );
  XOR2 MCInst1_MC1_v2_2Inst_1_U1  ( .A(MCInst1_MC1_v2_2Inst_1_n1 ), .B(
        MCInst1_MC1_v2_2Inst_1_n2 ), .Z(MCInst1_MC1_v2_2 [1]) );
  XOR2 MCInst1_MC1_v3_0Inst_1_U1  ( .A(MCInst1_MC1_v3_2 [2]), .B(
        MCInst1_MC1_v3_2 [3]), .Z(MCInst1_MC1_v3_0 [1]) );
  XOR2 MCInst1_MC1_v3_1Inst_1_U1  ( .A(MCInst1_MC1_v3_0 [3]), .B(
        MCInst1_MC1_v3_2 [3]), .Z(MCInst1_MC1_v3_1 [1]) );
  XOR2 MCInst1_MC1_v3_3Inst_1_U2  ( .A(MCInst1_MC1_v3_2 [2]), .B(
        MCInst1_MC1_v3_0 [3]), .Z(MCInst1_MC1_v3_3Inst_1_n1 ) );
  XOR2 MCInst1_MC1_v3_3Inst_1_U1  ( .A(MCInst1_MC1_v3_2 [3]), .B(
        MCInst1_MC1_v3_3Inst_1_n1 ), .Z(MCInst1_MC1_v3_3 [1]) );
  XOR2 MCInst1_MC1_v0_0Inst_2_U1  ( .A(MCInst1_MC1_v0_3 [0]), .B(
        ShiftRowsOutput[56]), .Z(MCInst1_MC1_v0_0 [2]) );
  XOR2 MCInst1_MC1_v0_1Inst_2_U1  ( .A(MCInst1_MC1_v0_3 [0]), .B(
        MCInst1_MC1_v0_3 [3]), .Z(MCInst1_MC1_v0_1 [2]) );
  XOR2 MCInst1_MC1_v0_2Inst_2_U1  ( .A(MCInst1_MC1_v0_3 [0]), .B(
        MCInst1_MC1_v0_0 [3]), .Z(MCInst1_MC1_v0_2 [2]) );
  XOR2 MCInst1_MC1_v1_1Inst_2_U2  ( .A(MCInst1_MC1_v1_3 [0]), .B(
        MCInst1_MC1_v1_3 [2]), .Z(MCInst1_MC1_v1_1Inst_2_n1 ) );
  XOR2 MCInst1_MC1_v1_1Inst_2_U1  ( .A(ShiftRowsOutput[40]), .B(
        MCInst1_MC1_v1_1Inst_2_n1 ), .Z(MCInst1_MC1_v1_1 [2]) );
  XOR2 MCInst1_MC1_v1_2Inst_2_U2  ( .A(MCInst1_MC1_v1_3 [3]), .B(
        MCInst1_MC1_v1_3 [2]), .Z(MCInst1_MC1_v1_2Inst_2_n1 ) );
  XOR2 MCInst1_MC1_v1_2Inst_2_U1  ( .A(ShiftRowsOutput[40]), .B(
        MCInst1_MC1_v1_2Inst_2_n1 ), .Z(MCInst1_MC1_v1_2 [2]) );
  XOR2 MCInst1_MC1_v2_1Inst_2_U2  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v2_0 [3]), .Z(MCInst1_MC1_v2_1Inst_2_n1 ) );
  XOR2 MCInst1_MC1_v2_1Inst_2_U1  ( .A(MCInst1_MC1_v2_3 [1]), .B(
        MCInst1_MC1_v2_1Inst_2_n1 ), .Z(MCInst1_MC1_v2_1 [2]) );
  XOR2 MCInst1_MC1_v2_2Inst_2_U2  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v2_0 [3]), .Z(MCInst1_MC1_v2_2Inst_2_n1 ) );
  XOR2 MCInst1_MC1_v2_2Inst_2_U1  ( .A(MCInst1_MC1_v2_0 [2]), .B(
        MCInst1_MC1_v2_2Inst_2_n1 ), .Z(MCInst1_MC1_v2_2 [2]) );
  XOR2 MCInst1_MC1_v2_3Inst_2_U1  ( .A(MCInst1_MC1_v2_0 [2]), .B(
        MCInst1_MC1_v2_3 [1]), .Z(MCInst1_MC1_v2_3 [2]) );
  XOR2 MCInst1_MC1_v3_1Inst_2_U2  ( .A(MCInst1_MC1_v3_2 [2]), .B(
        MCInst1_MC1_v3_0 [2]), .Z(MCInst1_MC1_v3_1Inst_2_n1 ) );
  XOR2 MCInst1_MC1_v3_1Inst_2_U1  ( .A(MCInst1_MC1_v3_2 [3]), .B(
        MCInst1_MC1_v3_1Inst_2_n1 ), .Z(MCInst1_MC1_v3_1 [2]) );
  XOR2 MCInst1_MC1_v3_3Inst_2_U1  ( .A(MCInst1_MC1_v3_2 [2]), .B(
        MCInst1_MC1_v3_0 [2]), .Z(MCInst1_MC1_v3_3 [2]) );
  XOR2 MCInst1_MC1_v0_1Inst_3_U1  ( .A(MCInst1_MC1_v0_3 [0]), .B(
        ShiftRowsOutput[56]), .Z(MCInst1_MC1_v0_1 [3]) );
  XOR2 MCInst1_MC1_v0_2Inst_3_U1  ( .A(MCInst1_MC1_v0_3 [3]), .B(
        ShiftRowsOutput[56]), .Z(MCInst1_MC1_v0_2 [3]) );
  XOR2 MCInst1_MC1_v1_1Inst_3_U1  ( .A(MCInst1_MC1_v1_3 [3]), .B(
        MCInst1_MC1_v1_3 [2]), .Z(MCInst1_MC1_v1_1 [3]) );
  XOR2 MCInst1_MC1_v1_2Inst_3_U3  ( .A(MCInst1_MC1_v1_3 [0]), .B(
        MCInst1_MC1_v1_3 [3]), .Z(MCInst1_MC1_v1_2Inst_3_n1 ) );
  XOR2 MCInst1_MC1_v1_2Inst_3_U2  ( .A(MCInst1_MC1_v1_3 [2]), .B(
        ShiftRowsOutput[40]), .Z(MCInst1_MC1_v1_2Inst_3_n2 ) );
  XOR2 MCInst1_MC1_v1_2Inst_3_U1  ( .A(MCInst1_MC1_v1_2Inst_3_n1 ), .B(
        MCInst1_MC1_v1_2Inst_3_n2 ), .Z(MCInst1_MC1_v1_2 [3]) );
  XOR2 MCInst1_MC1_v2_1Inst_3_U1  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v2_0 [2]), .Z(MCInst1_MC1_v2_1 [3]) );
  XOR2 MCInst1_MC1_v2_2Inst_3_U2  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v2_0 [3]), .Z(MCInst1_MC1_v2_2Inst_3_n1 ) );
  XOR2 MCInst1_MC1_v2_2Inst_3_U1  ( .A(MCInst1_MC1_v2_3 [1]), .B(
        MCInst1_MC1_v2_2Inst_3_n1 ), .Z(MCInst1_MC1_v2_2 [3]) );
  XOR2 MCInst1_MC1_v2_3Inst_3_U2  ( .A(MCInst1_MC1_v2_0 [3]), .B(
        MCInst1_MC1_v2_0 [2]), .Z(MCInst1_MC1_v2_3Inst_3_n1 ) );
  XOR2 MCInst1_MC1_v2_3Inst_3_U1  ( .A(MCInst1_MC1_v2_3 [1]), .B(
        MCInst1_MC1_v2_3Inst_3_n1 ), .Z(MCInst1_MC1_v2_3 [3]) );
  XOR2 MCInst1_MC1_v3_1Inst_3_U1  ( .A(MCInst1_MC1_v3_0 [3]), .B(
        MCInst1_MC1_v3_0 [2]), .Z(MCInst1_MC1_v3_1 [3]) );
  XOR2 MCInst1_MC1_v3_3Inst_3_U1  ( .A(MCInst1_MC1_v3_0 [3]), .B(
        MCInst1_MC1_v3_2 [3]), .Z(MCInst1_MC1_v3_3 [3]) );
  XOR2 MCInst1_MC1_r0Inst_XORInst_0_0_U4  ( .A(
        MCInst1_MC1_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC1_r0Inst_XORInst_0_0_n6 ), .Z(Feedback[56]) );
  XOR2 MCInst1_MC1_r0Inst_XORInst_0_0_U3  ( .A(1'b0), .B(
        MCInst1_MC1_r0Inst_XORInst_0_0_n4 ), .Z(
        MCInst1_MC1_r0Inst_XORInst_0_0_n6 ) );
  XOR2 MCInst1_MC1_r0Inst_XORInst_0_0_U2  ( .A(MCInst1_MC1_v2_0 [0]), .B(
        MCInst1_MC1_v3_2 [2]), .Z(MCInst1_MC1_r0Inst_XORInst_0_0_n5 ) );
  XOR2 MCInst1_MC1_r0Inst_XORInst_0_0_U1  ( .A(MCInst1_MC1_v0_3 [3]), .B(
        ShiftRowsOutput[40]), .Z(MCInst1_MC1_r0Inst_XORInst_0_0_n4 ) );
  XOR2 MCInst1_MC1_r0Inst_XORInst_0_1_U4  ( .A(
        MCInst1_MC1_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC1_r0Inst_XORInst_0_1_n6 ), .Z(Feedback[57]) );
  XOR2 MCInst1_MC1_r0Inst_XORInst_0_1_U3  ( .A(1'b0), .B(
        MCInst1_MC1_r0Inst_XORInst_0_1_n4 ), .Z(
        MCInst1_MC1_r0Inst_XORInst_0_1_n6 ) );
  XOR2 MCInst1_MC1_r0Inst_XORInst_0_1_U2  ( .A(MCInst1_MC1_v2_0 [1]), .B(
        MCInst1_MC1_v3_0 [1]), .Z(MCInst1_MC1_r0Inst_XORInst_0_1_n5 ) );
  XOR2 MCInst1_MC1_r0Inst_XORInst_0_1_U1  ( .A(MCInst1_MC1_v0_0 [1]), .B(
        MCInst1_MC1_v1_3 [2]), .Z(MCInst1_MC1_r0Inst_XORInst_0_1_n4 ) );
  XOR2 MCInst1_MC1_r0Inst_XORInst_0_2_U4  ( .A(
        MCInst1_MC1_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC1_r0Inst_XORInst_0_2_n6 ), .Z(Feedback[58]) );
  XOR2 MCInst1_MC1_r0Inst_XORInst_0_2_U3  ( .A(1'b0), .B(
        MCInst1_MC1_r0Inst_XORInst_0_2_n4 ), .Z(
        MCInst1_MC1_r0Inst_XORInst_0_2_n6 ) );
  XOR2 MCInst1_MC1_r0Inst_XORInst_0_2_U2  ( .A(MCInst1_MC1_v2_0 [2]), .B(
        MCInst1_MC1_v3_0 [2]), .Z(MCInst1_MC1_r0Inst_XORInst_0_2_n5 ) );
  XOR2 MCInst1_MC1_r0Inst_XORInst_0_2_U1  ( .A(MCInst1_MC1_v0_0 [2]), .B(
        MCInst1_MC1_v1_3 [3]), .Z(MCInst1_MC1_r0Inst_XORInst_0_2_n4 ) );
  XOR2 MCInst1_MC1_r0Inst_XORInst_0_3_U4  ( .A(
        MCInst1_MC1_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC1_r0Inst_XORInst_0_3_n6 ), .Z(Feedback[59]) );
  XOR2 MCInst1_MC1_r0Inst_XORInst_0_3_U3  ( .A(1'b0), .B(
        MCInst1_MC1_r0Inst_XORInst_0_3_n4 ), .Z(
        MCInst1_MC1_r0Inst_XORInst_0_3_n6 ) );
  XOR2 MCInst1_MC1_r0Inst_XORInst_0_3_U2  ( .A(MCInst1_MC1_v2_0 [3]), .B(
        MCInst1_MC1_v3_0 [3]), .Z(MCInst1_MC1_r0Inst_XORInst_0_3_n5 ) );
  XOR2 MCInst1_MC1_r0Inst_XORInst_0_3_U1  ( .A(MCInst1_MC1_v0_0 [3]), .B(
        MCInst1_MC1_v1_3 [0]), .Z(MCInst1_MC1_r0Inst_XORInst_0_3_n4 ) );
  XOR2 MCInst1_MC1_r1Inst_XORInst_0_0_U4  ( .A(
        MCInst1_MC1_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC1_r1Inst_XORInst_0_0_n6 ), .Z(Feedback[40]) );
  XOR2 MCInst1_MC1_r1Inst_XORInst_0_0_U3  ( .A(1'b0), .B(
        MCInst1_MC1_r1Inst_XORInst_0_0_n4 ), .Z(
        MCInst1_MC1_r1Inst_XORInst_0_0_n6 ) );
  XOR2 MCInst1_MC1_r1Inst_XORInst_0_0_U2  ( .A(MCInst1_MC1_v2_1 [0]), .B(
        MCInst1_MC1_v3_1 [0]), .Z(MCInst1_MC1_r1Inst_XORInst_0_0_n5 ) );
  XOR2 MCInst1_MC1_r1Inst_XORInst_0_0_U1  ( .A(MCInst1_MC1_v0_0 [3]), .B(
        MCInst1_MC1_v1_1 [0]), .Z(MCInst1_MC1_r1Inst_XORInst_0_0_n4 ) );
  XOR2 MCInst1_MC1_r1Inst_XORInst_0_1_U4  ( .A(
        MCInst1_MC1_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC1_r1Inst_XORInst_0_1_n6 ), .Z(Feedback[41]) );
  XOR2 MCInst1_MC1_r1Inst_XORInst_0_1_U3  ( .A(1'b0), .B(
        MCInst1_MC1_r1Inst_XORInst_0_1_n4 ), .Z(
        MCInst1_MC1_r1Inst_XORInst_0_1_n6 ) );
  XOR2 MCInst1_MC1_r1Inst_XORInst_0_1_U2  ( .A(MCInst1_MC1_v2_1 [1]), .B(
        MCInst1_MC1_v3_1 [1]), .Z(MCInst1_MC1_r1Inst_XORInst_0_1_n5 ) );
  XOR2 MCInst1_MC1_r1Inst_XORInst_0_1_U1  ( .A(MCInst1_MC1_v0_1 [1]), .B(
        MCInst1_MC1_v1_1 [1]), .Z(MCInst1_MC1_r1Inst_XORInst_0_1_n4 ) );
  XOR2 MCInst1_MC1_r1Inst_XORInst_0_2_U4  ( .A(
        MCInst1_MC1_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC1_r1Inst_XORInst_0_2_n6 ), .Z(Feedback[42]) );
  XOR2 MCInst1_MC1_r1Inst_XORInst_0_2_U3  ( .A(1'b0), .B(
        MCInst1_MC1_r1Inst_XORInst_0_2_n4 ), .Z(
        MCInst1_MC1_r1Inst_XORInst_0_2_n6 ) );
  XOR2 MCInst1_MC1_r1Inst_XORInst_0_2_U2  ( .A(MCInst1_MC1_v2_1 [2]), .B(
        MCInst1_MC1_v3_1 [2]), .Z(MCInst1_MC1_r1Inst_XORInst_0_2_n5 ) );
  XOR2 MCInst1_MC1_r1Inst_XORInst_0_2_U1  ( .A(MCInst1_MC1_v0_1 [2]), .B(
        MCInst1_MC1_v1_1 [2]), .Z(MCInst1_MC1_r1Inst_XORInst_0_2_n4 ) );
  XOR2 MCInst1_MC1_r1Inst_XORInst_0_3_U4  ( .A(
        MCInst1_MC1_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC1_r1Inst_XORInst_0_3_n6 ), .Z(Feedback[43]) );
  XOR2 MCInst1_MC1_r1Inst_XORInst_0_3_U3  ( .A(1'b0), .B(
        MCInst1_MC1_r1Inst_XORInst_0_3_n4 ), .Z(
        MCInst1_MC1_r1Inst_XORInst_0_3_n6 ) );
  XOR2 MCInst1_MC1_r1Inst_XORInst_0_3_U2  ( .A(MCInst1_MC1_v2_1 [3]), .B(
        MCInst1_MC1_v3_1 [3]), .Z(MCInst1_MC1_r1Inst_XORInst_0_3_n5 ) );
  XOR2 MCInst1_MC1_r1Inst_XORInst_0_3_U1  ( .A(MCInst1_MC1_v0_1 [3]), .B(
        MCInst1_MC1_v1_1 [3]), .Z(MCInst1_MC1_r1Inst_XORInst_0_3_n4 ) );
  XOR2 MCInst1_MC1_r2Inst_XORInst_0_0_U4  ( .A(
        MCInst1_MC1_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC1_r2Inst_XORInst_0_0_n6 ), .Z(Feedback[24]) );
  XOR2 MCInst1_MC1_r2Inst_XORInst_0_0_U3  ( .A(1'b0), .B(
        MCInst1_MC1_r2Inst_XORInst_0_0_n4 ), .Z(
        MCInst1_MC1_r2Inst_XORInst_0_0_n6 ) );
  XOR2 MCInst1_MC1_r2Inst_XORInst_0_0_U2  ( .A(MCInst1_MC1_v2_2 [0]), .B(
        MCInst1_MC1_v3_2 [0]), .Z(MCInst1_MC1_r2Inst_XORInst_0_0_n5 ) );
  XOR2 MCInst1_MC1_r2Inst_XORInst_0_0_U1  ( .A(MCInst1_MC1_v0_2 [0]), .B(
        MCInst1_MC1_v1_2 [0]), .Z(MCInst1_MC1_r2Inst_XORInst_0_0_n4 ) );
  XOR2 MCInst1_MC1_r2Inst_XORInst_0_1_U4  ( .A(
        MCInst1_MC1_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC1_r2Inst_XORInst_0_1_n6 ), .Z(Feedback[25]) );
  XOR2 MCInst1_MC1_r2Inst_XORInst_0_1_U3  ( .A(1'b0), .B(
        MCInst1_MC1_r2Inst_XORInst_0_1_n4 ), .Z(
        MCInst1_MC1_r2Inst_XORInst_0_1_n6 ) );
  XOR2 MCInst1_MC1_r2Inst_XORInst_0_1_U2  ( .A(MCInst1_MC1_v2_2 [1]), .B(
        MCInst1_MC1_v3_0 [3]), .Z(MCInst1_MC1_r2Inst_XORInst_0_1_n5 ) );
  XOR2 MCInst1_MC1_r2Inst_XORInst_0_1_U1  ( .A(MCInst1_MC1_v0_2 [1]), .B(
        MCInst1_MC1_v1_2 [1]), .Z(MCInst1_MC1_r2Inst_XORInst_0_1_n4 ) );
  XOR2 MCInst1_MC1_r2Inst_XORInst_0_2_U4  ( .A(
        MCInst1_MC1_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC1_r2Inst_XORInst_0_2_n6 ), .Z(Feedback[26]) );
  XOR2 MCInst1_MC1_r2Inst_XORInst_0_2_U3  ( .A(1'b0), .B(
        MCInst1_MC1_r2Inst_XORInst_0_2_n4 ), .Z(
        MCInst1_MC1_r2Inst_XORInst_0_2_n6 ) );
  XOR2 MCInst1_MC1_r2Inst_XORInst_0_2_U2  ( .A(MCInst1_MC1_v2_2 [2]), .B(
        MCInst1_MC1_v3_2 [2]), .Z(MCInst1_MC1_r2Inst_XORInst_0_2_n5 ) );
  XOR2 MCInst1_MC1_r2Inst_XORInst_0_2_U1  ( .A(MCInst1_MC1_v0_2 [2]), .B(
        MCInst1_MC1_v1_2 [2]), .Z(MCInst1_MC1_r2Inst_XORInst_0_2_n4 ) );
  XOR2 MCInst1_MC1_r2Inst_XORInst_0_3_U4  ( .A(
        MCInst1_MC1_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC1_r2Inst_XORInst_0_3_n6 ), .Z(Feedback[27]) );
  XOR2 MCInst1_MC1_r2Inst_XORInst_0_3_U3  ( .A(1'b0), .B(
        MCInst1_MC1_r2Inst_XORInst_0_3_n4 ), .Z(
        MCInst1_MC1_r2Inst_XORInst_0_3_n6 ) );
  XOR2 MCInst1_MC1_r2Inst_XORInst_0_3_U2  ( .A(MCInst1_MC1_v2_2 [3]), .B(
        MCInst1_MC1_v3_2 [3]), .Z(MCInst1_MC1_r2Inst_XORInst_0_3_n5 ) );
  XOR2 MCInst1_MC1_r2Inst_XORInst_0_3_U1  ( .A(MCInst1_MC1_v0_2 [3]), .B(
        MCInst1_MC1_v1_2 [3]), .Z(MCInst1_MC1_r2Inst_XORInst_0_3_n4 ) );
  XOR2 MCInst1_MC1_r3Inst_XORInst_0_0_U4  ( .A(
        MCInst1_MC1_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC1_r3Inst_XORInst_0_0_n6 ), .Z(Feedback[8]) );
  XOR2 MCInst1_MC1_r3Inst_XORInst_0_0_U3  ( .A(1'b0), .B(
        MCInst1_MC1_r3Inst_XORInst_0_0_n4 ), .Z(
        MCInst1_MC1_r3Inst_XORInst_0_0_n6 ) );
  XOR2 MCInst1_MC1_r3Inst_XORInst_0_0_U2  ( .A(MCInst1_MC1_v2_3 [0]), .B(
        MCInst1_MC1_v3_3 [0]), .Z(MCInst1_MC1_r3Inst_XORInst_0_0_n5 ) );
  XOR2 MCInst1_MC1_r3Inst_XORInst_0_0_U1  ( .A(MCInst1_MC1_v0_3 [0]), .B(
        MCInst1_MC1_v1_3 [0]), .Z(MCInst1_MC1_r3Inst_XORInst_0_0_n4 ) );
  XOR2 MCInst1_MC1_r3Inst_XORInst_0_1_U4  ( .A(
        MCInst1_MC1_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC1_r3Inst_XORInst_0_1_n6 ), .Z(Feedback[9]) );
  XOR2 MCInst1_MC1_r3Inst_XORInst_0_1_U3  ( .A(1'b0), .B(
        MCInst1_MC1_r3Inst_XORInst_0_1_n4 ), .Z(
        MCInst1_MC1_r3Inst_XORInst_0_1_n6 ) );
  XOR2 MCInst1_MC1_r3Inst_XORInst_0_1_U2  ( .A(MCInst1_MC1_v2_3 [1]), .B(
        MCInst1_MC1_v3_3 [1]), .Z(MCInst1_MC1_r3Inst_XORInst_0_1_n5 ) );
  XOR2 MCInst1_MC1_r3Inst_XORInst_0_1_U1  ( .A(MCInst1_MC1_v0_3 [1]), .B(
        MCInst1_MC1_v1_3 [1]), .Z(MCInst1_MC1_r3Inst_XORInst_0_1_n4 ) );
  XOR2 MCInst1_MC1_r3Inst_XORInst_0_2_U4  ( .A(
        MCInst1_MC1_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC1_r3Inst_XORInst_0_2_n6 ), .Z(Feedback[10]) );
  XOR2 MCInst1_MC1_r3Inst_XORInst_0_2_U3  ( .A(1'b0), .B(
        MCInst1_MC1_r3Inst_XORInst_0_2_n4 ), .Z(
        MCInst1_MC1_r3Inst_XORInst_0_2_n6 ) );
  XOR2 MCInst1_MC1_r3Inst_XORInst_0_2_U2  ( .A(MCInst1_MC1_v2_3 [2]), .B(
        MCInst1_MC1_v3_3 [2]), .Z(MCInst1_MC1_r3Inst_XORInst_0_2_n5 ) );
  XOR2 MCInst1_MC1_r3Inst_XORInst_0_2_U1  ( .A(MCInst1_MC1_v0_0 [3]), .B(
        MCInst1_MC1_v1_3 [2]), .Z(MCInst1_MC1_r3Inst_XORInst_0_2_n4 ) );
  XOR2 MCInst1_MC1_r3Inst_XORInst_0_3_U4  ( .A(
        MCInst1_MC1_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC1_r3Inst_XORInst_0_3_n6 ), .Z(Feedback[11]) );
  XOR2 MCInst1_MC1_r3Inst_XORInst_0_3_U3  ( .A(1'b0), .B(
        MCInst1_MC1_r3Inst_XORInst_0_3_n4 ), .Z(
        MCInst1_MC1_r3Inst_XORInst_0_3_n6 ) );
  XOR2 MCInst1_MC1_r3Inst_XORInst_0_3_U2  ( .A(MCInst1_MC1_v2_3 [3]), .B(
        MCInst1_MC1_v3_3 [3]), .Z(MCInst1_MC1_r3Inst_XORInst_0_3_n5 ) );
  XOR2 MCInst1_MC1_r3Inst_XORInst_0_3_U1  ( .A(MCInst1_MC1_v0_3 [3]), .B(
        MCInst1_MC1_v1_3 [3]), .Z(MCInst1_MC1_r3Inst_XORInst_0_3_n4 ) );
  XOR2 MCInst1_MC2_v0_2Inst_0_U2  ( .A(MCInst1_MC2_v0_3 [0]), .B(
        MCInst1_MC2_v0_0 [3]), .Z(MCInst1_MC2_v0_2Inst_0_n1 ) );
  XOR2 MCInst1_MC2_v0_2Inst_0_U1  ( .A(ShiftRowsOutput[52]), .B(
        MCInst1_MC2_v0_2Inst_0_n1 ), .Z(MCInst1_MC2_v0_2 [0]) );
  XOR2 MCInst1_MC2_v1_1Inst_0_U1  ( .A(MCInst1_MC2_v1_3 [0]), .B(
        MCInst1_MC2_v1_3 [3]), .Z(MCInst1_MC2_v1_1 [0]) );
  XOR2 MCInst1_MC2_v1_2Inst_0_U2  ( .A(MCInst1_MC2_v1_3 [0]), .B(
        MCInst1_MC2_v1_3 [3]), .Z(MCInst1_MC2_v1_2Inst_0_n1 ) );
  XOR2 MCInst1_MC2_v1_2Inst_0_U1  ( .A(MCInst1_MC2_v1_3 [2]), .B(
        MCInst1_MC2_v1_2Inst_0_n1 ), .Z(MCInst1_MC2_v1_2 [0]) );
  XOR2 MCInst1_MC2_v2_1Inst_0_U1  ( .A(MCInst1_MC2_v2_0 [3]), .B(
        MCInst1_MC2_v2_3 [1]), .Z(MCInst1_MC2_v2_1 [0]) );
  XOR2 MCInst1_MC2_v2_2Inst_0_U1  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v2_0 [2]), .Z(MCInst1_MC2_v2_2 [0]) );
  XOR2 MCInst1_MC2_v2_3Inst_0_U3  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v2_0 [3]), .Z(MCInst1_MC2_v2_3Inst_0_n1 ) );
  XOR2 MCInst1_MC2_v2_3Inst_0_U2  ( .A(MCInst1_MC2_v2_0 [2]), .B(
        MCInst1_MC2_v2_3 [1]), .Z(MCInst1_MC2_v2_3Inst_0_n2 ) );
  XOR2 MCInst1_MC2_v2_3Inst_0_U1  ( .A(MCInst1_MC2_v2_3Inst_0_n1 ), .B(
        MCInst1_MC2_v2_3Inst_0_n2 ), .Z(MCInst1_MC2_v2_3 [0]) );
  XOR2 MCInst1_MC2_v3_1Inst_0_U1  ( .A(MCInst1_MC2_v3_2 [2]), .B(
        MCInst1_MC2_v3_0 [3]), .Z(MCInst1_MC2_v3_1 [0]) );
  XOR2 MCInst1_MC2_v3_2Inst_0_U1  ( .A(MCInst1_MC2_v3_0 [2]), .B(
        MCInst1_MC2_v3_2 [3]), .Z(MCInst1_MC2_v3_2 [0]) );
  XOR2 MCInst1_MC2_v3_3Inst_0_U2  ( .A(MCInst1_MC2_v3_2 [2]), .B(
        MCInst1_MC2_v3_0 [2]), .Z(MCInst1_MC2_v3_3Inst_0_n1 ) );
  XOR2 MCInst1_MC2_v3_3Inst_0_U1  ( .A(MCInst1_MC2_v3_2 [3]), .B(
        MCInst1_MC2_v3_3Inst_0_n1 ), .Z(MCInst1_MC2_v3_3 [0]) );
  XOR2 MCInst1_MC2_v0_0Inst_1_U1  ( .A(MCInst1_MC2_v0_3 [0]), .B(
        MCInst1_MC2_v0_3 [3]), .Z(MCInst1_MC2_v0_0 [1]) );
  XOR2 MCInst1_MC2_v0_1Inst_1_U1  ( .A(MCInst1_MC2_v0_3 [3]), .B(
        MCInst1_MC2_v0_0 [3]), .Z(MCInst1_MC2_v0_1 [1]) );
  XOR2 MCInst1_MC2_v0_2Inst_1_U2  ( .A(MCInst1_MC2_v0_3 [0]), .B(
        MCInst1_MC2_v0_3 [3]), .Z(MCInst1_MC2_v0_2Inst_1_n1 ) );
  XOR2 MCInst1_MC2_v0_2Inst_1_U1  ( .A(ShiftRowsOutput[52]), .B(
        MCInst1_MC2_v0_2Inst_1_n1 ), .Z(MCInst1_MC2_v0_2 [1]) );
  XOR2 MCInst1_MC2_v0_3Inst_1_U1  ( .A(MCInst1_MC2_v0_3 [0]), .B(
        ShiftRowsOutput[52]), .Z(MCInst1_MC2_v0_3 [1]) );
  XOR2 MCInst1_MC2_v1_1Inst_1_U1  ( .A(MCInst1_MC2_v1_3 [3]), .B(
        ShiftRowsOutput[36]), .Z(MCInst1_MC2_v1_1 [1]) );
  XOR2 MCInst1_MC2_v1_2Inst_1_U1  ( .A(MCInst1_MC2_v1_3 [2]), .B(
        ShiftRowsOutput[36]), .Z(MCInst1_MC2_v1_2 [1]) );
  XOR2 MCInst1_MC2_v1_3Inst_1_U1  ( .A(MCInst1_MC2_v1_3 [0]), .B(
        ShiftRowsOutput[36]), .Z(MCInst1_MC2_v1_3 [1]) );
  XOR2 MCInst1_MC2_v2_0Inst_1_U1  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v2_3 [1]), .Z(MCInst1_MC2_v2_0 [1]) );
  XOR2 MCInst1_MC2_v2_1Inst_1_U2  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v2_0 [3]), .Z(MCInst1_MC2_v2_1Inst_1_n1 ) );
  XOR2 MCInst1_MC2_v2_1Inst_1_U1  ( .A(MCInst1_MC2_v2_0 [2]), .B(
        MCInst1_MC2_v2_1Inst_1_n1 ), .Z(MCInst1_MC2_v2_1 [1]) );
  XOR2 MCInst1_MC2_v2_2Inst_1_U3  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v2_0 [3]), .Z(MCInst1_MC2_v2_2Inst_1_n1 ) );
  XOR2 MCInst1_MC2_v2_2Inst_1_U2  ( .A(MCInst1_MC2_v2_0 [2]), .B(
        MCInst1_MC2_v2_3 [1]), .Z(MCInst1_MC2_v2_2Inst_1_n2 ) );
  XOR2 MCInst1_MC2_v2_2Inst_1_U1  ( .A(MCInst1_MC2_v2_2Inst_1_n1 ), .B(
        MCInst1_MC2_v2_2Inst_1_n2 ), .Z(MCInst1_MC2_v2_2 [1]) );
  XOR2 MCInst1_MC2_v3_0Inst_1_U1  ( .A(MCInst1_MC2_v3_2 [2]), .B(
        MCInst1_MC2_v3_2 [3]), .Z(MCInst1_MC2_v3_0 [1]) );
  XOR2 MCInst1_MC2_v3_1Inst_1_U1  ( .A(MCInst1_MC2_v3_0 [3]), .B(
        MCInst1_MC2_v3_2 [3]), .Z(MCInst1_MC2_v3_1 [1]) );
  XOR2 MCInst1_MC2_v3_3Inst_1_U2  ( .A(MCInst1_MC2_v3_2 [2]), .B(
        MCInst1_MC2_v3_0 [3]), .Z(MCInst1_MC2_v3_3Inst_1_n1 ) );
  XOR2 MCInst1_MC2_v3_3Inst_1_U1  ( .A(MCInst1_MC2_v3_2 [3]), .B(
        MCInst1_MC2_v3_3Inst_1_n1 ), .Z(MCInst1_MC2_v3_3 [1]) );
  XOR2 MCInst1_MC2_v0_0Inst_2_U1  ( .A(MCInst1_MC2_v0_3 [0]), .B(
        ShiftRowsOutput[52]), .Z(MCInst1_MC2_v0_0 [2]) );
  XOR2 MCInst1_MC2_v0_1Inst_2_U1  ( .A(MCInst1_MC2_v0_3 [0]), .B(
        MCInst1_MC2_v0_3 [3]), .Z(MCInst1_MC2_v0_1 [2]) );
  XOR2 MCInst1_MC2_v0_2Inst_2_U1  ( .A(MCInst1_MC2_v0_3 [0]), .B(
        MCInst1_MC2_v0_0 [3]), .Z(MCInst1_MC2_v0_2 [2]) );
  XOR2 MCInst1_MC2_v1_1Inst_2_U2  ( .A(MCInst1_MC2_v1_3 [0]), .B(
        MCInst1_MC2_v1_3 [2]), .Z(MCInst1_MC2_v1_1Inst_2_n1 ) );
  XOR2 MCInst1_MC2_v1_1Inst_2_U1  ( .A(ShiftRowsOutput[36]), .B(
        MCInst1_MC2_v1_1Inst_2_n1 ), .Z(MCInst1_MC2_v1_1 [2]) );
  XOR2 MCInst1_MC2_v1_2Inst_2_U2  ( .A(MCInst1_MC2_v1_3 [3]), .B(
        MCInst1_MC2_v1_3 [2]), .Z(MCInst1_MC2_v1_2Inst_2_n1 ) );
  XOR2 MCInst1_MC2_v1_2Inst_2_U1  ( .A(ShiftRowsOutput[36]), .B(
        MCInst1_MC2_v1_2Inst_2_n1 ), .Z(MCInst1_MC2_v1_2 [2]) );
  XOR2 MCInst1_MC2_v2_1Inst_2_U2  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v2_0 [3]), .Z(MCInst1_MC2_v2_1Inst_2_n1 ) );
  XOR2 MCInst1_MC2_v2_1Inst_2_U1  ( .A(MCInst1_MC2_v2_3 [1]), .B(
        MCInst1_MC2_v2_1Inst_2_n1 ), .Z(MCInst1_MC2_v2_1 [2]) );
  XOR2 MCInst1_MC2_v2_2Inst_2_U2  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v2_0 [3]), .Z(MCInst1_MC2_v2_2Inst_2_n1 ) );
  XOR2 MCInst1_MC2_v2_2Inst_2_U1  ( .A(MCInst1_MC2_v2_0 [2]), .B(
        MCInst1_MC2_v2_2Inst_2_n1 ), .Z(MCInst1_MC2_v2_2 [2]) );
  XOR2 MCInst1_MC2_v2_3Inst_2_U1  ( .A(MCInst1_MC2_v2_0 [2]), .B(
        MCInst1_MC2_v2_3 [1]), .Z(MCInst1_MC2_v2_3 [2]) );
  XOR2 MCInst1_MC2_v3_1Inst_2_U2  ( .A(MCInst1_MC2_v3_2 [2]), .B(
        MCInst1_MC2_v3_0 [2]), .Z(MCInst1_MC2_v3_1Inst_2_n1 ) );
  XOR2 MCInst1_MC2_v3_1Inst_2_U1  ( .A(MCInst1_MC2_v3_2 [3]), .B(
        MCInst1_MC2_v3_1Inst_2_n1 ), .Z(MCInst1_MC2_v3_1 [2]) );
  XOR2 MCInst1_MC2_v3_3Inst_2_U1  ( .A(MCInst1_MC2_v3_2 [2]), .B(
        MCInst1_MC2_v3_0 [2]), .Z(MCInst1_MC2_v3_3 [2]) );
  XOR2 MCInst1_MC2_v0_1Inst_3_U1  ( .A(MCInst1_MC2_v0_3 [0]), .B(
        ShiftRowsOutput[52]), .Z(MCInst1_MC2_v0_1 [3]) );
  XOR2 MCInst1_MC2_v0_2Inst_3_U1  ( .A(MCInst1_MC2_v0_3 [3]), .B(
        ShiftRowsOutput[52]), .Z(MCInst1_MC2_v0_2 [3]) );
  XOR2 MCInst1_MC2_v1_1Inst_3_U1  ( .A(MCInst1_MC2_v1_3 [3]), .B(
        MCInst1_MC2_v1_3 [2]), .Z(MCInst1_MC2_v1_1 [3]) );
  XOR2 MCInst1_MC2_v1_2Inst_3_U3  ( .A(MCInst1_MC2_v1_3 [0]), .B(
        MCInst1_MC2_v1_3 [3]), .Z(MCInst1_MC2_v1_2Inst_3_n1 ) );
  XOR2 MCInst1_MC2_v1_2Inst_3_U2  ( .A(MCInst1_MC2_v1_3 [2]), .B(
        ShiftRowsOutput[36]), .Z(MCInst1_MC2_v1_2Inst_3_n2 ) );
  XOR2 MCInst1_MC2_v1_2Inst_3_U1  ( .A(MCInst1_MC2_v1_2Inst_3_n1 ), .B(
        MCInst1_MC2_v1_2Inst_3_n2 ), .Z(MCInst1_MC2_v1_2 [3]) );
  XOR2 MCInst1_MC2_v2_1Inst_3_U1  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v2_0 [2]), .Z(MCInst1_MC2_v2_1 [3]) );
  XOR2 MCInst1_MC2_v2_2Inst_3_U2  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v2_0 [3]), .Z(MCInst1_MC2_v2_2Inst_3_n1 ) );
  XOR2 MCInst1_MC2_v2_2Inst_3_U1  ( .A(MCInst1_MC2_v2_3 [1]), .B(
        MCInst1_MC2_v2_2Inst_3_n1 ), .Z(MCInst1_MC2_v2_2 [3]) );
  XOR2 MCInst1_MC2_v2_3Inst_3_U2  ( .A(MCInst1_MC2_v2_0 [3]), .B(
        MCInst1_MC2_v2_0 [2]), .Z(MCInst1_MC2_v2_3Inst_3_n1 ) );
  XOR2 MCInst1_MC2_v2_3Inst_3_U1  ( .A(MCInst1_MC2_v2_3 [1]), .B(
        MCInst1_MC2_v2_3Inst_3_n1 ), .Z(MCInst1_MC2_v2_3 [3]) );
  XOR2 MCInst1_MC2_v3_1Inst_3_U1  ( .A(MCInst1_MC2_v3_0 [3]), .B(
        MCInst1_MC2_v3_0 [2]), .Z(MCInst1_MC2_v3_1 [3]) );
  XOR2 MCInst1_MC2_v3_3Inst_3_U1  ( .A(MCInst1_MC2_v3_0 [3]), .B(
        MCInst1_MC2_v3_2 [3]), .Z(MCInst1_MC2_v3_3 [3]) );
  XOR2 MCInst1_MC2_r0Inst_XORInst_0_0_U4  ( .A(
        MCInst1_MC2_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC2_r0Inst_XORInst_0_0_n6 ), .Z(Feedback[52]) );
  XOR2 MCInst1_MC2_r0Inst_XORInst_0_0_U3  ( .A(1'b0), .B(
        MCInst1_MC2_r0Inst_XORInst_0_0_n4 ), .Z(
        MCInst1_MC2_r0Inst_XORInst_0_0_n6 ) );
  XOR2 MCInst1_MC2_r0Inst_XORInst_0_0_U2  ( .A(MCInst1_MC2_v2_0 [0]), .B(
        MCInst1_MC2_v3_2 [2]), .Z(MCInst1_MC2_r0Inst_XORInst_0_0_n5 ) );
  XOR2 MCInst1_MC2_r0Inst_XORInst_0_0_U1  ( .A(MCInst1_MC2_v0_3 [3]), .B(
        ShiftRowsOutput[36]), .Z(MCInst1_MC2_r0Inst_XORInst_0_0_n4 ) );
  XOR2 MCInst1_MC2_r0Inst_XORInst_0_1_U4  ( .A(
        MCInst1_MC2_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC2_r0Inst_XORInst_0_1_n6 ), .Z(Feedback[53]) );
  XOR2 MCInst1_MC2_r0Inst_XORInst_0_1_U3  ( .A(1'b0), .B(
        MCInst1_MC2_r0Inst_XORInst_0_1_n4 ), .Z(
        MCInst1_MC2_r0Inst_XORInst_0_1_n6 ) );
  XOR2 MCInst1_MC2_r0Inst_XORInst_0_1_U2  ( .A(MCInst1_MC2_v2_0 [1]), .B(
        MCInst1_MC2_v3_0 [1]), .Z(MCInst1_MC2_r0Inst_XORInst_0_1_n5 ) );
  XOR2 MCInst1_MC2_r0Inst_XORInst_0_1_U1  ( .A(MCInst1_MC2_v0_0 [1]), .B(
        MCInst1_MC2_v1_3 [2]), .Z(MCInst1_MC2_r0Inst_XORInst_0_1_n4 ) );
  XOR2 MCInst1_MC2_r0Inst_XORInst_0_2_U4  ( .A(
        MCInst1_MC2_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC2_r0Inst_XORInst_0_2_n6 ), .Z(Feedback[54]) );
  XOR2 MCInst1_MC2_r0Inst_XORInst_0_2_U3  ( .A(1'b0), .B(
        MCInst1_MC2_r0Inst_XORInst_0_2_n4 ), .Z(
        MCInst1_MC2_r0Inst_XORInst_0_2_n6 ) );
  XOR2 MCInst1_MC2_r0Inst_XORInst_0_2_U2  ( .A(MCInst1_MC2_v2_0 [2]), .B(
        MCInst1_MC2_v3_0 [2]), .Z(MCInst1_MC2_r0Inst_XORInst_0_2_n5 ) );
  XOR2 MCInst1_MC2_r0Inst_XORInst_0_2_U1  ( .A(MCInst1_MC2_v0_0 [2]), .B(
        MCInst1_MC2_v1_3 [3]), .Z(MCInst1_MC2_r0Inst_XORInst_0_2_n4 ) );
  XOR2 MCInst1_MC2_r0Inst_XORInst_0_3_U4  ( .A(
        MCInst1_MC2_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC2_r0Inst_XORInst_0_3_n6 ), .Z(Feedback[55]) );
  XOR2 MCInst1_MC2_r0Inst_XORInst_0_3_U3  ( .A(1'b0), .B(
        MCInst1_MC2_r0Inst_XORInst_0_3_n4 ), .Z(
        MCInst1_MC2_r0Inst_XORInst_0_3_n6 ) );
  XOR2 MCInst1_MC2_r0Inst_XORInst_0_3_U2  ( .A(MCInst1_MC2_v2_0 [3]), .B(
        MCInst1_MC2_v3_0 [3]), .Z(MCInst1_MC2_r0Inst_XORInst_0_3_n5 ) );
  XOR2 MCInst1_MC2_r0Inst_XORInst_0_3_U1  ( .A(MCInst1_MC2_v0_0 [3]), .B(
        MCInst1_MC2_v1_3 [0]), .Z(MCInst1_MC2_r0Inst_XORInst_0_3_n4 ) );
  XOR2 MCInst1_MC2_r1Inst_XORInst_0_0_U4  ( .A(
        MCInst1_MC2_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC2_r1Inst_XORInst_0_0_n6 ), .Z(Feedback[36]) );
  XOR2 MCInst1_MC2_r1Inst_XORInst_0_0_U3  ( .A(1'b0), .B(
        MCInst1_MC2_r1Inst_XORInst_0_0_n4 ), .Z(
        MCInst1_MC2_r1Inst_XORInst_0_0_n6 ) );
  XOR2 MCInst1_MC2_r1Inst_XORInst_0_0_U2  ( .A(MCInst1_MC2_v2_1 [0]), .B(
        MCInst1_MC2_v3_1 [0]), .Z(MCInst1_MC2_r1Inst_XORInst_0_0_n5 ) );
  XOR2 MCInst1_MC2_r1Inst_XORInst_0_0_U1  ( .A(MCInst1_MC2_v0_0 [3]), .B(
        MCInst1_MC2_v1_1 [0]), .Z(MCInst1_MC2_r1Inst_XORInst_0_0_n4 ) );
  XOR2 MCInst1_MC2_r1Inst_XORInst_0_1_U4  ( .A(
        MCInst1_MC2_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC2_r1Inst_XORInst_0_1_n6 ), .Z(Feedback[37]) );
  XOR2 MCInst1_MC2_r1Inst_XORInst_0_1_U3  ( .A(1'b0), .B(
        MCInst1_MC2_r1Inst_XORInst_0_1_n4 ), .Z(
        MCInst1_MC2_r1Inst_XORInst_0_1_n6 ) );
  XOR2 MCInst1_MC2_r1Inst_XORInst_0_1_U2  ( .A(MCInst1_MC2_v2_1 [1]), .B(
        MCInst1_MC2_v3_1 [1]), .Z(MCInst1_MC2_r1Inst_XORInst_0_1_n5 ) );
  XOR2 MCInst1_MC2_r1Inst_XORInst_0_1_U1  ( .A(MCInst1_MC2_v0_1 [1]), .B(
        MCInst1_MC2_v1_1 [1]), .Z(MCInst1_MC2_r1Inst_XORInst_0_1_n4 ) );
  XOR2 MCInst1_MC2_r1Inst_XORInst_0_2_U4  ( .A(
        MCInst1_MC2_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC2_r1Inst_XORInst_0_2_n6 ), .Z(Feedback[38]) );
  XOR2 MCInst1_MC2_r1Inst_XORInst_0_2_U3  ( .A(1'b0), .B(
        MCInst1_MC2_r1Inst_XORInst_0_2_n4 ), .Z(
        MCInst1_MC2_r1Inst_XORInst_0_2_n6 ) );
  XOR2 MCInst1_MC2_r1Inst_XORInst_0_2_U2  ( .A(MCInst1_MC2_v2_1 [2]), .B(
        MCInst1_MC2_v3_1 [2]), .Z(MCInst1_MC2_r1Inst_XORInst_0_2_n5 ) );
  XOR2 MCInst1_MC2_r1Inst_XORInst_0_2_U1  ( .A(MCInst1_MC2_v0_1 [2]), .B(
        MCInst1_MC2_v1_1 [2]), .Z(MCInst1_MC2_r1Inst_XORInst_0_2_n4 ) );
  XOR2 MCInst1_MC2_r1Inst_XORInst_0_3_U4  ( .A(
        MCInst1_MC2_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC2_r1Inst_XORInst_0_3_n6 ), .Z(Feedback[39]) );
  XOR2 MCInst1_MC2_r1Inst_XORInst_0_3_U3  ( .A(1'b0), .B(
        MCInst1_MC2_r1Inst_XORInst_0_3_n4 ), .Z(
        MCInst1_MC2_r1Inst_XORInst_0_3_n6 ) );
  XOR2 MCInst1_MC2_r1Inst_XORInst_0_3_U2  ( .A(MCInst1_MC2_v2_1 [3]), .B(
        MCInst1_MC2_v3_1 [3]), .Z(MCInst1_MC2_r1Inst_XORInst_0_3_n5 ) );
  XOR2 MCInst1_MC2_r1Inst_XORInst_0_3_U1  ( .A(MCInst1_MC2_v0_1 [3]), .B(
        MCInst1_MC2_v1_1 [3]), .Z(MCInst1_MC2_r1Inst_XORInst_0_3_n4 ) );
  XOR2 MCInst1_MC2_r2Inst_XORInst_0_0_U4  ( .A(
        MCInst1_MC2_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC2_r2Inst_XORInst_0_0_n6 ), .Z(Feedback[20]) );
  XOR2 MCInst1_MC2_r2Inst_XORInst_0_0_U3  ( .A(1'b0), .B(
        MCInst1_MC2_r2Inst_XORInst_0_0_n4 ), .Z(
        MCInst1_MC2_r2Inst_XORInst_0_0_n6 ) );
  XOR2 MCInst1_MC2_r2Inst_XORInst_0_0_U2  ( .A(MCInst1_MC2_v2_2 [0]), .B(
        MCInst1_MC2_v3_2 [0]), .Z(MCInst1_MC2_r2Inst_XORInst_0_0_n5 ) );
  XOR2 MCInst1_MC2_r2Inst_XORInst_0_0_U1  ( .A(MCInst1_MC2_v0_2 [0]), .B(
        MCInst1_MC2_v1_2 [0]), .Z(MCInst1_MC2_r2Inst_XORInst_0_0_n4 ) );
  XOR2 MCInst1_MC2_r2Inst_XORInst_0_1_U4  ( .A(
        MCInst1_MC2_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC2_r2Inst_XORInst_0_1_n6 ), .Z(Feedback[21]) );
  XOR2 MCInst1_MC2_r2Inst_XORInst_0_1_U3  ( .A(1'b0), .B(
        MCInst1_MC2_r2Inst_XORInst_0_1_n4 ), .Z(
        MCInst1_MC2_r2Inst_XORInst_0_1_n6 ) );
  XOR2 MCInst1_MC2_r2Inst_XORInst_0_1_U2  ( .A(MCInst1_MC2_v2_2 [1]), .B(
        MCInst1_MC2_v3_0 [3]), .Z(MCInst1_MC2_r2Inst_XORInst_0_1_n5 ) );
  XOR2 MCInst1_MC2_r2Inst_XORInst_0_1_U1  ( .A(MCInst1_MC2_v0_2 [1]), .B(
        MCInst1_MC2_v1_2 [1]), .Z(MCInst1_MC2_r2Inst_XORInst_0_1_n4 ) );
  XOR2 MCInst1_MC2_r2Inst_XORInst_0_2_U4  ( .A(
        MCInst1_MC2_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC2_r2Inst_XORInst_0_2_n6 ), .Z(Feedback[22]) );
  XOR2 MCInst1_MC2_r2Inst_XORInst_0_2_U3  ( .A(1'b0), .B(
        MCInst1_MC2_r2Inst_XORInst_0_2_n4 ), .Z(
        MCInst1_MC2_r2Inst_XORInst_0_2_n6 ) );
  XOR2 MCInst1_MC2_r2Inst_XORInst_0_2_U2  ( .A(MCInst1_MC2_v2_2 [2]), .B(
        MCInst1_MC2_v3_2 [2]), .Z(MCInst1_MC2_r2Inst_XORInst_0_2_n5 ) );
  XOR2 MCInst1_MC2_r2Inst_XORInst_0_2_U1  ( .A(MCInst1_MC2_v0_2 [2]), .B(
        MCInst1_MC2_v1_2 [2]), .Z(MCInst1_MC2_r2Inst_XORInst_0_2_n4 ) );
  XOR2 MCInst1_MC2_r2Inst_XORInst_0_3_U4  ( .A(
        MCInst1_MC2_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC2_r2Inst_XORInst_0_3_n6 ), .Z(Feedback[23]) );
  XOR2 MCInst1_MC2_r2Inst_XORInst_0_3_U3  ( .A(1'b0), .B(
        MCInst1_MC2_r2Inst_XORInst_0_3_n4 ), .Z(
        MCInst1_MC2_r2Inst_XORInst_0_3_n6 ) );
  XOR2 MCInst1_MC2_r2Inst_XORInst_0_3_U2  ( .A(MCInst1_MC2_v2_2 [3]), .B(
        MCInst1_MC2_v3_2 [3]), .Z(MCInst1_MC2_r2Inst_XORInst_0_3_n5 ) );
  XOR2 MCInst1_MC2_r2Inst_XORInst_0_3_U1  ( .A(MCInst1_MC2_v0_2 [3]), .B(
        MCInst1_MC2_v1_2 [3]), .Z(MCInst1_MC2_r2Inst_XORInst_0_3_n4 ) );
  XOR2 MCInst1_MC2_r3Inst_XORInst_0_0_U4  ( .A(
        MCInst1_MC2_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC2_r3Inst_XORInst_0_0_n6 ), .Z(Feedback[4]) );
  XOR2 MCInst1_MC2_r3Inst_XORInst_0_0_U3  ( .A(1'b0), .B(
        MCInst1_MC2_r3Inst_XORInst_0_0_n4 ), .Z(
        MCInst1_MC2_r3Inst_XORInst_0_0_n6 ) );
  XOR2 MCInst1_MC2_r3Inst_XORInst_0_0_U2  ( .A(MCInst1_MC2_v2_3 [0]), .B(
        MCInst1_MC2_v3_3 [0]), .Z(MCInst1_MC2_r3Inst_XORInst_0_0_n5 ) );
  XOR2 MCInst1_MC2_r3Inst_XORInst_0_0_U1  ( .A(MCInst1_MC2_v0_3 [0]), .B(
        MCInst1_MC2_v1_3 [0]), .Z(MCInst1_MC2_r3Inst_XORInst_0_0_n4 ) );
  XOR2 MCInst1_MC2_r3Inst_XORInst_0_1_U4  ( .A(
        MCInst1_MC2_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC2_r3Inst_XORInst_0_1_n6 ), .Z(Feedback[5]) );
  XOR2 MCInst1_MC2_r3Inst_XORInst_0_1_U3  ( .A(1'b0), .B(
        MCInst1_MC2_r3Inst_XORInst_0_1_n4 ), .Z(
        MCInst1_MC2_r3Inst_XORInst_0_1_n6 ) );
  XOR2 MCInst1_MC2_r3Inst_XORInst_0_1_U2  ( .A(MCInst1_MC2_v2_3 [1]), .B(
        MCInst1_MC2_v3_3 [1]), .Z(MCInst1_MC2_r3Inst_XORInst_0_1_n5 ) );
  XOR2 MCInst1_MC2_r3Inst_XORInst_0_1_U1  ( .A(MCInst1_MC2_v0_3 [1]), .B(
        MCInst1_MC2_v1_3 [1]), .Z(MCInst1_MC2_r3Inst_XORInst_0_1_n4 ) );
  XOR2 MCInst1_MC2_r3Inst_XORInst_0_2_U4  ( .A(
        MCInst1_MC2_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC2_r3Inst_XORInst_0_2_n6 ), .Z(Feedback[6]) );
  XOR2 MCInst1_MC2_r3Inst_XORInst_0_2_U3  ( .A(1'b0), .B(
        MCInst1_MC2_r3Inst_XORInst_0_2_n4 ), .Z(
        MCInst1_MC2_r3Inst_XORInst_0_2_n6 ) );
  XOR2 MCInst1_MC2_r3Inst_XORInst_0_2_U2  ( .A(MCInst1_MC2_v2_3 [2]), .B(
        MCInst1_MC2_v3_3 [2]), .Z(MCInst1_MC2_r3Inst_XORInst_0_2_n5 ) );
  XOR2 MCInst1_MC2_r3Inst_XORInst_0_2_U1  ( .A(MCInst1_MC2_v0_0 [3]), .B(
        MCInst1_MC2_v1_3 [2]), .Z(MCInst1_MC2_r3Inst_XORInst_0_2_n4 ) );
  XOR2 MCInst1_MC2_r3Inst_XORInst_0_3_U4  ( .A(
        MCInst1_MC2_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC2_r3Inst_XORInst_0_3_n6 ), .Z(Feedback[7]) );
  XOR2 MCInst1_MC2_r3Inst_XORInst_0_3_U3  ( .A(1'b0), .B(
        MCInst1_MC2_r3Inst_XORInst_0_3_n4 ), .Z(
        MCInst1_MC2_r3Inst_XORInst_0_3_n6 ) );
  XOR2 MCInst1_MC2_r3Inst_XORInst_0_3_U2  ( .A(MCInst1_MC2_v2_3 [3]), .B(
        MCInst1_MC2_v3_3 [3]), .Z(MCInst1_MC2_r3Inst_XORInst_0_3_n5 ) );
  XOR2 MCInst1_MC2_r3Inst_XORInst_0_3_U1  ( .A(MCInst1_MC2_v0_3 [3]), .B(
        MCInst1_MC2_v1_3 [3]), .Z(MCInst1_MC2_r3Inst_XORInst_0_3_n4 ) );
  XOR2 MCInst1_MC3_v0_2Inst_0_U2  ( .A(MCInst1_MC3_v0_3 [0]), .B(
        MCInst1_MC3_v0_0 [3]), .Z(MCInst1_MC3_v0_2Inst_0_n1 ) );
  XOR2 MCInst1_MC3_v0_2Inst_0_U1  ( .A(ShiftRowsOutput[48]), .B(
        MCInst1_MC3_v0_2Inst_0_n1 ), .Z(MCInst1_MC3_v0_2 [0]) );
  XOR2 MCInst1_MC3_v1_1Inst_0_U1  ( .A(MCInst1_MC3_v1_3 [0]), .B(
        MCInst1_MC3_v1_3 [3]), .Z(MCInst1_MC3_v1_1 [0]) );
  XOR2 MCInst1_MC3_v1_2Inst_0_U2  ( .A(MCInst1_MC3_v1_3 [0]), .B(
        MCInst1_MC3_v1_3 [3]), .Z(MCInst1_MC3_v1_2Inst_0_n1 ) );
  XOR2 MCInst1_MC3_v1_2Inst_0_U1  ( .A(MCInst1_MC3_v1_3 [2]), .B(
        MCInst1_MC3_v1_2Inst_0_n1 ), .Z(MCInst1_MC3_v1_2 [0]) );
  XOR2 MCInst1_MC3_v2_1Inst_0_U1  ( .A(MCInst1_MC3_v2_0 [3]), .B(
        MCInst1_MC3_v2_3 [1]), .Z(MCInst1_MC3_v2_1 [0]) );
  XOR2 MCInst1_MC3_v2_2Inst_0_U1  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v2_0 [2]), .Z(MCInst1_MC3_v2_2 [0]) );
  XOR2 MCInst1_MC3_v2_3Inst_0_U3  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v2_0 [3]), .Z(MCInst1_MC3_v2_3Inst_0_n1 ) );
  XOR2 MCInst1_MC3_v2_3Inst_0_U2  ( .A(MCInst1_MC3_v2_0 [2]), .B(
        MCInst1_MC3_v2_3 [1]), .Z(MCInst1_MC3_v2_3Inst_0_n2 ) );
  XOR2 MCInst1_MC3_v2_3Inst_0_U1  ( .A(MCInst1_MC3_v2_3Inst_0_n1 ), .B(
        MCInst1_MC3_v2_3Inst_0_n2 ), .Z(MCInst1_MC3_v2_3 [0]) );
  XOR2 MCInst1_MC3_v3_1Inst_0_U1  ( .A(MCInst1_MC3_v3_2 [2]), .B(
        MCInst1_MC3_v3_0 [3]), .Z(MCInst1_MC3_v3_1 [0]) );
  XOR2 MCInst1_MC3_v3_2Inst_0_U1  ( .A(MCInst1_MC3_v3_0 [2]), .B(
        MCInst1_MC3_v3_2 [3]), .Z(MCInst1_MC3_v3_2 [0]) );
  XOR2 MCInst1_MC3_v3_3Inst_0_U2  ( .A(MCInst1_MC3_v3_2 [2]), .B(
        MCInst1_MC3_v3_0 [2]), .Z(MCInst1_MC3_v3_3Inst_0_n1 ) );
  XOR2 MCInst1_MC3_v3_3Inst_0_U1  ( .A(MCInst1_MC3_v3_2 [3]), .B(
        MCInst1_MC3_v3_3Inst_0_n1 ), .Z(MCInst1_MC3_v3_3 [0]) );
  XOR2 MCInst1_MC3_v0_0Inst_1_U1  ( .A(MCInst1_MC3_v0_3 [0]), .B(
        MCInst1_MC3_v0_3 [3]), .Z(MCInst1_MC3_v0_0 [1]) );
  XOR2 MCInst1_MC3_v0_1Inst_1_U1  ( .A(MCInst1_MC3_v0_3 [3]), .B(
        MCInst1_MC3_v0_0 [3]), .Z(MCInst1_MC3_v0_1 [1]) );
  XOR2 MCInst1_MC3_v0_2Inst_1_U2  ( .A(MCInst1_MC3_v0_3 [0]), .B(
        MCInst1_MC3_v0_3 [3]), .Z(MCInst1_MC3_v0_2Inst_1_n1 ) );
  XOR2 MCInst1_MC3_v0_2Inst_1_U1  ( .A(ShiftRowsOutput[48]), .B(
        MCInst1_MC3_v0_2Inst_1_n1 ), .Z(MCInst1_MC3_v0_2 [1]) );
  XOR2 MCInst1_MC3_v0_3Inst_1_U1  ( .A(MCInst1_MC3_v0_3 [0]), .B(
        ShiftRowsOutput[48]), .Z(MCInst1_MC3_v0_3 [1]) );
  XOR2 MCInst1_MC3_v1_1Inst_1_U1  ( .A(MCInst1_MC3_v1_3 [3]), .B(
        ShiftRowsOutput[32]), .Z(MCInst1_MC3_v1_1 [1]) );
  XOR2 MCInst1_MC3_v1_2Inst_1_U1  ( .A(MCInst1_MC3_v1_3 [2]), .B(
        ShiftRowsOutput[32]), .Z(MCInst1_MC3_v1_2 [1]) );
  XOR2 MCInst1_MC3_v1_3Inst_1_U1  ( .A(MCInst1_MC3_v1_3 [0]), .B(
        ShiftRowsOutput[32]), .Z(MCInst1_MC3_v1_3 [1]) );
  XOR2 MCInst1_MC3_v2_0Inst_1_U1  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v2_3 [1]), .Z(MCInst1_MC3_v2_0 [1]) );
  XOR2 MCInst1_MC3_v2_1Inst_1_U2  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v2_0 [3]), .Z(MCInst1_MC3_v2_1Inst_1_n1 ) );
  XOR2 MCInst1_MC3_v2_1Inst_1_U1  ( .A(MCInst1_MC3_v2_0 [2]), .B(
        MCInst1_MC3_v2_1Inst_1_n1 ), .Z(MCInst1_MC3_v2_1 [1]) );
  XOR2 MCInst1_MC3_v2_2Inst_1_U3  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v2_0 [3]), .Z(MCInst1_MC3_v2_2Inst_1_n1 ) );
  XOR2 MCInst1_MC3_v2_2Inst_1_U2  ( .A(MCInst1_MC3_v2_0 [2]), .B(
        MCInst1_MC3_v2_3 [1]), .Z(MCInst1_MC3_v2_2Inst_1_n2 ) );
  XOR2 MCInst1_MC3_v2_2Inst_1_U1  ( .A(MCInst1_MC3_v2_2Inst_1_n1 ), .B(
        MCInst1_MC3_v2_2Inst_1_n2 ), .Z(MCInst1_MC3_v2_2 [1]) );
  XOR2 MCInst1_MC3_v3_0Inst_1_U1  ( .A(MCInst1_MC3_v3_2 [2]), .B(
        MCInst1_MC3_v3_2 [3]), .Z(MCInst1_MC3_v3_0 [1]) );
  XOR2 MCInst1_MC3_v3_1Inst_1_U1  ( .A(MCInst1_MC3_v3_0 [3]), .B(
        MCInst1_MC3_v3_2 [3]), .Z(MCInst1_MC3_v3_1 [1]) );
  XOR2 MCInst1_MC3_v3_3Inst_1_U2  ( .A(MCInst1_MC3_v3_2 [2]), .B(
        MCInst1_MC3_v3_0 [3]), .Z(MCInst1_MC3_v3_3Inst_1_n1 ) );
  XOR2 MCInst1_MC3_v3_3Inst_1_U1  ( .A(MCInst1_MC3_v3_2 [3]), .B(
        MCInst1_MC3_v3_3Inst_1_n1 ), .Z(MCInst1_MC3_v3_3 [1]) );
  XOR2 MCInst1_MC3_v0_0Inst_2_U1  ( .A(MCInst1_MC3_v0_3 [0]), .B(
        ShiftRowsOutput[48]), .Z(MCInst1_MC3_v0_0 [2]) );
  XOR2 MCInst1_MC3_v0_1Inst_2_U1  ( .A(MCInst1_MC3_v0_3 [0]), .B(
        MCInst1_MC3_v0_3 [3]), .Z(MCInst1_MC3_v0_1 [2]) );
  XOR2 MCInst1_MC3_v0_2Inst_2_U1  ( .A(MCInst1_MC3_v0_3 [0]), .B(
        MCInst1_MC3_v0_0 [3]), .Z(MCInst1_MC3_v0_2 [2]) );
  XOR2 MCInst1_MC3_v1_1Inst_2_U2  ( .A(MCInst1_MC3_v1_3 [0]), .B(
        MCInst1_MC3_v1_3 [2]), .Z(MCInst1_MC3_v1_1Inst_2_n1 ) );
  XOR2 MCInst1_MC3_v1_1Inst_2_U1  ( .A(ShiftRowsOutput[32]), .B(
        MCInst1_MC3_v1_1Inst_2_n1 ), .Z(MCInst1_MC3_v1_1 [2]) );
  XOR2 MCInst1_MC3_v1_2Inst_2_U2  ( .A(MCInst1_MC3_v1_3 [3]), .B(
        MCInst1_MC3_v1_3 [2]), .Z(MCInst1_MC3_v1_2Inst_2_n1 ) );
  XOR2 MCInst1_MC3_v1_2Inst_2_U1  ( .A(ShiftRowsOutput[32]), .B(
        MCInst1_MC3_v1_2Inst_2_n1 ), .Z(MCInst1_MC3_v1_2 [2]) );
  XOR2 MCInst1_MC3_v2_1Inst_2_U2  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v2_0 [3]), .Z(MCInst1_MC3_v2_1Inst_2_n1 ) );
  XOR2 MCInst1_MC3_v2_1Inst_2_U1  ( .A(MCInst1_MC3_v2_3 [1]), .B(
        MCInst1_MC3_v2_1Inst_2_n1 ), .Z(MCInst1_MC3_v2_1 [2]) );
  XOR2 MCInst1_MC3_v2_2Inst_2_U2  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v2_0 [3]), .Z(MCInst1_MC3_v2_2Inst_2_n1 ) );
  XOR2 MCInst1_MC3_v2_2Inst_2_U1  ( .A(MCInst1_MC3_v2_0 [2]), .B(
        MCInst1_MC3_v2_2Inst_2_n1 ), .Z(MCInst1_MC3_v2_2 [2]) );
  XOR2 MCInst1_MC3_v2_3Inst_2_U1  ( .A(MCInst1_MC3_v2_0 [2]), .B(
        MCInst1_MC3_v2_3 [1]), .Z(MCInst1_MC3_v2_3 [2]) );
  XOR2 MCInst1_MC3_v3_1Inst_2_U2  ( .A(MCInst1_MC3_v3_2 [2]), .B(
        MCInst1_MC3_v3_0 [2]), .Z(MCInst1_MC3_v3_1Inst_2_n1 ) );
  XOR2 MCInst1_MC3_v3_1Inst_2_U1  ( .A(MCInst1_MC3_v3_2 [3]), .B(
        MCInst1_MC3_v3_1Inst_2_n1 ), .Z(MCInst1_MC3_v3_1 [2]) );
  XOR2 MCInst1_MC3_v3_3Inst_2_U1  ( .A(MCInst1_MC3_v3_2 [2]), .B(
        MCInst1_MC3_v3_0 [2]), .Z(MCInst1_MC3_v3_3 [2]) );
  XOR2 MCInst1_MC3_v0_1Inst_3_U1  ( .A(MCInst1_MC3_v0_3 [0]), .B(
        ShiftRowsOutput[48]), .Z(MCInst1_MC3_v0_1 [3]) );
  XOR2 MCInst1_MC3_v0_2Inst_3_U1  ( .A(MCInst1_MC3_v0_3 [3]), .B(
        ShiftRowsOutput[48]), .Z(MCInst1_MC3_v0_2 [3]) );
  XOR2 MCInst1_MC3_v1_1Inst_3_U1  ( .A(MCInst1_MC3_v1_3 [3]), .B(
        MCInst1_MC3_v1_3 [2]), .Z(MCInst1_MC3_v1_1 [3]) );
  XOR2 MCInst1_MC3_v1_2Inst_3_U3  ( .A(MCInst1_MC3_v1_3 [0]), .B(
        MCInst1_MC3_v1_3 [3]), .Z(MCInst1_MC3_v1_2Inst_3_n1 ) );
  XOR2 MCInst1_MC3_v1_2Inst_3_U2  ( .A(MCInst1_MC3_v1_3 [2]), .B(
        ShiftRowsOutput[32]), .Z(MCInst1_MC3_v1_2Inst_3_n2 ) );
  XOR2 MCInst1_MC3_v1_2Inst_3_U1  ( .A(MCInst1_MC3_v1_2Inst_3_n1 ), .B(
        MCInst1_MC3_v1_2Inst_3_n2 ), .Z(MCInst1_MC3_v1_2 [3]) );
  XOR2 MCInst1_MC3_v2_1Inst_3_U1  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v2_0 [2]), .Z(MCInst1_MC3_v2_1 [3]) );
  XOR2 MCInst1_MC3_v2_2Inst_3_U2  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v2_0 [3]), .Z(MCInst1_MC3_v2_2Inst_3_n1 ) );
  XOR2 MCInst1_MC3_v2_2Inst_3_U1  ( .A(MCInst1_MC3_v2_3 [1]), .B(
        MCInst1_MC3_v2_2Inst_3_n1 ), .Z(MCInst1_MC3_v2_2 [3]) );
  XOR2 MCInst1_MC3_v2_3Inst_3_U2  ( .A(MCInst1_MC3_v2_0 [3]), .B(
        MCInst1_MC3_v2_0 [2]), .Z(MCInst1_MC3_v2_3Inst_3_n1 ) );
  XOR2 MCInst1_MC3_v2_3Inst_3_U1  ( .A(MCInst1_MC3_v2_3 [1]), .B(
        MCInst1_MC3_v2_3Inst_3_n1 ), .Z(MCInst1_MC3_v2_3 [3]) );
  XOR2 MCInst1_MC3_v3_1Inst_3_U1  ( .A(MCInst1_MC3_v3_0 [3]), .B(
        MCInst1_MC3_v3_0 [2]), .Z(MCInst1_MC3_v3_1 [3]) );
  XOR2 MCInst1_MC3_v3_3Inst_3_U1  ( .A(MCInst1_MC3_v3_0 [3]), .B(
        MCInst1_MC3_v3_2 [3]), .Z(MCInst1_MC3_v3_3 [3]) );
  XOR2 MCInst1_MC3_r0Inst_XORInst_0_0_U4  ( .A(
        MCInst1_MC3_r0Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC3_r0Inst_XORInst_0_0_n6 ), .Z(Feedback[48]) );
  XOR2 MCInst1_MC3_r0Inst_XORInst_0_0_U3  ( .A(1'b0), .B(
        MCInst1_MC3_r0Inst_XORInst_0_0_n4 ), .Z(
        MCInst1_MC3_r0Inst_XORInst_0_0_n6 ) );
  XOR2 MCInst1_MC3_r0Inst_XORInst_0_0_U2  ( .A(MCInst1_MC3_v2_0 [0]), .B(
        MCInst1_MC3_v3_2 [2]), .Z(MCInst1_MC3_r0Inst_XORInst_0_0_n5 ) );
  XOR2 MCInst1_MC3_r0Inst_XORInst_0_0_U1  ( .A(MCInst1_MC3_v0_3 [3]), .B(
        ShiftRowsOutput[32]), .Z(MCInst1_MC3_r0Inst_XORInst_0_0_n4 ) );
  XOR2 MCInst1_MC3_r0Inst_XORInst_0_1_U4  ( .A(
        MCInst1_MC3_r0Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC3_r0Inst_XORInst_0_1_n6 ), .Z(Feedback[49]) );
  XOR2 MCInst1_MC3_r0Inst_XORInst_0_1_U3  ( .A(1'b0), .B(
        MCInst1_MC3_r0Inst_XORInst_0_1_n4 ), .Z(
        MCInst1_MC3_r0Inst_XORInst_0_1_n6 ) );
  XOR2 MCInst1_MC3_r0Inst_XORInst_0_1_U2  ( .A(MCInst1_MC3_v2_0 [1]), .B(
        MCInst1_MC3_v3_0 [1]), .Z(MCInst1_MC3_r0Inst_XORInst_0_1_n5 ) );
  XOR2 MCInst1_MC3_r0Inst_XORInst_0_1_U1  ( .A(MCInst1_MC3_v0_0 [1]), .B(
        MCInst1_MC3_v1_3 [2]), .Z(MCInst1_MC3_r0Inst_XORInst_0_1_n4 ) );
  XOR2 MCInst1_MC3_r0Inst_XORInst_0_2_U4  ( .A(
        MCInst1_MC3_r0Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC3_r0Inst_XORInst_0_2_n6 ), .Z(Feedback[50]) );
  XOR2 MCInst1_MC3_r0Inst_XORInst_0_2_U3  ( .A(1'b0), .B(
        MCInst1_MC3_r0Inst_XORInst_0_2_n4 ), .Z(
        MCInst1_MC3_r0Inst_XORInst_0_2_n6 ) );
  XOR2 MCInst1_MC3_r0Inst_XORInst_0_2_U2  ( .A(MCInst1_MC3_v2_0 [2]), .B(
        MCInst1_MC3_v3_0 [2]), .Z(MCInst1_MC3_r0Inst_XORInst_0_2_n5 ) );
  XOR2 MCInst1_MC3_r0Inst_XORInst_0_2_U1  ( .A(MCInst1_MC3_v0_0 [2]), .B(
        MCInst1_MC3_v1_3 [3]), .Z(MCInst1_MC3_r0Inst_XORInst_0_2_n4 ) );
  XOR2 MCInst1_MC3_r0Inst_XORInst_0_3_U4  ( .A(
        MCInst1_MC3_r0Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC3_r0Inst_XORInst_0_3_n6 ), .Z(Feedback[51]) );
  XOR2 MCInst1_MC3_r0Inst_XORInst_0_3_U3  ( .A(1'b0), .B(
        MCInst1_MC3_r0Inst_XORInst_0_3_n4 ), .Z(
        MCInst1_MC3_r0Inst_XORInst_0_3_n6 ) );
  XOR2 MCInst1_MC3_r0Inst_XORInst_0_3_U2  ( .A(MCInst1_MC3_v2_0 [3]), .B(
        MCInst1_MC3_v3_0 [3]), .Z(MCInst1_MC3_r0Inst_XORInst_0_3_n5 ) );
  XOR2 MCInst1_MC3_r0Inst_XORInst_0_3_U1  ( .A(MCInst1_MC3_v0_0 [3]), .B(
        MCInst1_MC3_v1_3 [0]), .Z(MCInst1_MC3_r0Inst_XORInst_0_3_n4 ) );
  XOR2 MCInst1_MC3_r1Inst_XORInst_0_0_U4  ( .A(
        MCInst1_MC3_r1Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC3_r1Inst_XORInst_0_0_n6 ), .Z(Feedback[32]) );
  XOR2 MCInst1_MC3_r1Inst_XORInst_0_0_U3  ( .A(1'b0), .B(
        MCInst1_MC3_r1Inst_XORInst_0_0_n4 ), .Z(
        MCInst1_MC3_r1Inst_XORInst_0_0_n6 ) );
  XOR2 MCInst1_MC3_r1Inst_XORInst_0_0_U2  ( .A(MCInst1_MC3_v2_1 [0]), .B(
        MCInst1_MC3_v3_1 [0]), .Z(MCInst1_MC3_r1Inst_XORInst_0_0_n5 ) );
  XOR2 MCInst1_MC3_r1Inst_XORInst_0_0_U1  ( .A(MCInst1_MC3_v0_0 [3]), .B(
        MCInst1_MC3_v1_1 [0]), .Z(MCInst1_MC3_r1Inst_XORInst_0_0_n4 ) );
  XOR2 MCInst1_MC3_r1Inst_XORInst_0_1_U4  ( .A(
        MCInst1_MC3_r1Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC3_r1Inst_XORInst_0_1_n6 ), .Z(Feedback[33]) );
  XOR2 MCInst1_MC3_r1Inst_XORInst_0_1_U3  ( .A(1'b0), .B(
        MCInst1_MC3_r1Inst_XORInst_0_1_n4 ), .Z(
        MCInst1_MC3_r1Inst_XORInst_0_1_n6 ) );
  XOR2 MCInst1_MC3_r1Inst_XORInst_0_1_U2  ( .A(MCInst1_MC3_v2_1 [1]), .B(
        MCInst1_MC3_v3_1 [1]), .Z(MCInst1_MC3_r1Inst_XORInst_0_1_n5 ) );
  XOR2 MCInst1_MC3_r1Inst_XORInst_0_1_U1  ( .A(MCInst1_MC3_v0_1 [1]), .B(
        MCInst1_MC3_v1_1 [1]), .Z(MCInst1_MC3_r1Inst_XORInst_0_1_n4 ) );
  XOR2 MCInst1_MC3_r1Inst_XORInst_0_2_U4  ( .A(
        MCInst1_MC3_r1Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC3_r1Inst_XORInst_0_2_n6 ), .Z(Feedback[34]) );
  XOR2 MCInst1_MC3_r1Inst_XORInst_0_2_U3  ( .A(1'b0), .B(
        MCInst1_MC3_r1Inst_XORInst_0_2_n4 ), .Z(
        MCInst1_MC3_r1Inst_XORInst_0_2_n6 ) );
  XOR2 MCInst1_MC3_r1Inst_XORInst_0_2_U2  ( .A(MCInst1_MC3_v2_1 [2]), .B(
        MCInst1_MC3_v3_1 [2]), .Z(MCInst1_MC3_r1Inst_XORInst_0_2_n5 ) );
  XOR2 MCInst1_MC3_r1Inst_XORInst_0_2_U1  ( .A(MCInst1_MC3_v0_1 [2]), .B(
        MCInst1_MC3_v1_1 [2]), .Z(MCInst1_MC3_r1Inst_XORInst_0_2_n4 ) );
  XOR2 MCInst1_MC3_r1Inst_XORInst_0_3_U4  ( .A(
        MCInst1_MC3_r1Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC3_r1Inst_XORInst_0_3_n6 ), .Z(Feedback[35]) );
  XOR2 MCInst1_MC3_r1Inst_XORInst_0_3_U3  ( .A(1'b0), .B(
        MCInst1_MC3_r1Inst_XORInst_0_3_n4 ), .Z(
        MCInst1_MC3_r1Inst_XORInst_0_3_n6 ) );
  XOR2 MCInst1_MC3_r1Inst_XORInst_0_3_U2  ( .A(MCInst1_MC3_v2_1 [3]), .B(
        MCInst1_MC3_v3_1 [3]), .Z(MCInst1_MC3_r1Inst_XORInst_0_3_n5 ) );
  XOR2 MCInst1_MC3_r1Inst_XORInst_0_3_U1  ( .A(MCInst1_MC3_v0_1 [3]), .B(
        MCInst1_MC3_v1_1 [3]), .Z(MCInst1_MC3_r1Inst_XORInst_0_3_n4 ) );
  XOR2 MCInst1_MC3_r2Inst_XORInst_0_0_U4  ( .A(
        MCInst1_MC3_r2Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC3_r2Inst_XORInst_0_0_n6 ), .Z(Feedback[16]) );
  XOR2 MCInst1_MC3_r2Inst_XORInst_0_0_U3  ( .A(1'b0), .B(
        MCInst1_MC3_r2Inst_XORInst_0_0_n4 ), .Z(
        MCInst1_MC3_r2Inst_XORInst_0_0_n6 ) );
  XOR2 MCInst1_MC3_r2Inst_XORInst_0_0_U2  ( .A(MCInst1_MC3_v2_2 [0]), .B(
        MCInst1_MC3_v3_2 [0]), .Z(MCInst1_MC3_r2Inst_XORInst_0_0_n5 ) );
  XOR2 MCInst1_MC3_r2Inst_XORInst_0_0_U1  ( .A(MCInst1_MC3_v0_2 [0]), .B(
        MCInst1_MC3_v1_2 [0]), .Z(MCInst1_MC3_r2Inst_XORInst_0_0_n4 ) );
  XOR2 MCInst1_MC3_r2Inst_XORInst_0_1_U4  ( .A(
        MCInst1_MC3_r2Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC3_r2Inst_XORInst_0_1_n6 ), .Z(Feedback[17]) );
  XOR2 MCInst1_MC3_r2Inst_XORInst_0_1_U3  ( .A(1'b0), .B(
        MCInst1_MC3_r2Inst_XORInst_0_1_n4 ), .Z(
        MCInst1_MC3_r2Inst_XORInst_0_1_n6 ) );
  XOR2 MCInst1_MC3_r2Inst_XORInst_0_1_U2  ( .A(MCInst1_MC3_v2_2 [1]), .B(
        MCInst1_MC3_v3_0 [3]), .Z(MCInst1_MC3_r2Inst_XORInst_0_1_n5 ) );
  XOR2 MCInst1_MC3_r2Inst_XORInst_0_1_U1  ( .A(MCInst1_MC3_v0_2 [1]), .B(
        MCInst1_MC3_v1_2 [1]), .Z(MCInst1_MC3_r2Inst_XORInst_0_1_n4 ) );
  XOR2 MCInst1_MC3_r2Inst_XORInst_0_2_U4  ( .A(
        MCInst1_MC3_r2Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC3_r2Inst_XORInst_0_2_n6 ), .Z(Feedback[18]) );
  XOR2 MCInst1_MC3_r2Inst_XORInst_0_2_U3  ( .A(1'b0), .B(
        MCInst1_MC3_r2Inst_XORInst_0_2_n4 ), .Z(
        MCInst1_MC3_r2Inst_XORInst_0_2_n6 ) );
  XOR2 MCInst1_MC3_r2Inst_XORInst_0_2_U2  ( .A(MCInst1_MC3_v2_2 [2]), .B(
        MCInst1_MC3_v3_2 [2]), .Z(MCInst1_MC3_r2Inst_XORInst_0_2_n5 ) );
  XOR2 MCInst1_MC3_r2Inst_XORInst_0_2_U1  ( .A(MCInst1_MC3_v0_2 [2]), .B(
        MCInst1_MC3_v1_2 [2]), .Z(MCInst1_MC3_r2Inst_XORInst_0_2_n4 ) );
  XOR2 MCInst1_MC3_r2Inst_XORInst_0_3_U4  ( .A(
        MCInst1_MC3_r2Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC3_r2Inst_XORInst_0_3_n6 ), .Z(Feedback[19]) );
  XOR2 MCInst1_MC3_r2Inst_XORInst_0_3_U3  ( .A(1'b0), .B(
        MCInst1_MC3_r2Inst_XORInst_0_3_n4 ), .Z(
        MCInst1_MC3_r2Inst_XORInst_0_3_n6 ) );
  XOR2 MCInst1_MC3_r2Inst_XORInst_0_3_U2  ( .A(MCInst1_MC3_v2_2 [3]), .B(
        MCInst1_MC3_v3_2 [3]), .Z(MCInst1_MC3_r2Inst_XORInst_0_3_n5 ) );
  XOR2 MCInst1_MC3_r2Inst_XORInst_0_3_U1  ( .A(MCInst1_MC3_v0_2 [3]), .B(
        MCInst1_MC3_v1_2 [3]), .Z(MCInst1_MC3_r2Inst_XORInst_0_3_n4 ) );
  XOR2 MCInst1_MC3_r3Inst_XORInst_0_0_U4  ( .A(
        MCInst1_MC3_r3Inst_XORInst_0_0_n5 ), .B(
        MCInst1_MC3_r3Inst_XORInst_0_0_n6 ), .Z(Feedback[0]) );
  XOR2 MCInst1_MC3_r3Inst_XORInst_0_0_U3  ( .A(1'b0), .B(
        MCInst1_MC3_r3Inst_XORInst_0_0_n4 ), .Z(
        MCInst1_MC3_r3Inst_XORInst_0_0_n6 ) );
  XOR2 MCInst1_MC3_r3Inst_XORInst_0_0_U2  ( .A(MCInst1_MC3_v2_3 [0]), .B(
        MCInst1_MC3_v3_3 [0]), .Z(MCInst1_MC3_r3Inst_XORInst_0_0_n5 ) );
  XOR2 MCInst1_MC3_r3Inst_XORInst_0_0_U1  ( .A(MCInst1_MC3_v0_3 [0]), .B(
        MCInst1_MC3_v1_3 [0]), .Z(MCInst1_MC3_r3Inst_XORInst_0_0_n4 ) );
  XOR2 MCInst1_MC3_r3Inst_XORInst_0_1_U4  ( .A(
        MCInst1_MC3_r3Inst_XORInst_0_1_n5 ), .B(
        MCInst1_MC3_r3Inst_XORInst_0_1_n6 ), .Z(Feedback[1]) );
  XOR2 MCInst1_MC3_r3Inst_XORInst_0_1_U3  ( .A(1'b0), .B(
        MCInst1_MC3_r3Inst_XORInst_0_1_n4 ), .Z(
        MCInst1_MC3_r3Inst_XORInst_0_1_n6 ) );
  XOR2 MCInst1_MC3_r3Inst_XORInst_0_1_U2  ( .A(MCInst1_MC3_v2_3 [1]), .B(
        MCInst1_MC3_v3_3 [1]), .Z(MCInst1_MC3_r3Inst_XORInst_0_1_n5 ) );
  XOR2 MCInst1_MC3_r3Inst_XORInst_0_1_U1  ( .A(MCInst1_MC3_v0_3 [1]), .B(
        MCInst1_MC3_v1_3 [1]), .Z(MCInst1_MC3_r3Inst_XORInst_0_1_n4 ) );
  XOR2 MCInst1_MC3_r3Inst_XORInst_0_2_U4  ( .A(
        MCInst1_MC3_r3Inst_XORInst_0_2_n5 ), .B(
        MCInst1_MC3_r3Inst_XORInst_0_2_n6 ), .Z(Feedback[2]) );
  XOR2 MCInst1_MC3_r3Inst_XORInst_0_2_U3  ( .A(1'b0), .B(
        MCInst1_MC3_r3Inst_XORInst_0_2_n4 ), .Z(
        MCInst1_MC3_r3Inst_XORInst_0_2_n6 ) );
  XOR2 MCInst1_MC3_r3Inst_XORInst_0_2_U2  ( .A(MCInst1_MC3_v2_3 [2]), .B(
        MCInst1_MC3_v3_3 [2]), .Z(MCInst1_MC3_r3Inst_XORInst_0_2_n5 ) );
  XOR2 MCInst1_MC3_r3Inst_XORInst_0_2_U1  ( .A(MCInst1_MC3_v0_0 [3]), .B(
        MCInst1_MC3_v1_3 [2]), .Z(MCInst1_MC3_r3Inst_XORInst_0_2_n4 ) );
  XOR2 MCInst1_MC3_r3Inst_XORInst_0_3_U4  ( .A(
        MCInst1_MC3_r3Inst_XORInst_0_3_n5 ), .B(
        MCInst1_MC3_r3Inst_XORInst_0_3_n6 ), .Z(Feedback[3]) );
  XOR2 MCInst1_MC3_r3Inst_XORInst_0_3_U3  ( .A(1'b0), .B(
        MCInst1_MC3_r3Inst_XORInst_0_3_n4 ), .Z(
        MCInst1_MC3_r3Inst_XORInst_0_3_n6 ) );
  XOR2 MCInst1_MC3_r3Inst_XORInst_0_3_U2  ( .A(MCInst1_MC3_v2_3 [3]), .B(
        MCInst1_MC3_v3_3 [3]), .Z(MCInst1_MC3_r3Inst_XORInst_0_3_n5 ) );
  XOR2 MCInst1_MC3_r3Inst_XORInst_0_3_U1  ( .A(MCInst1_MC3_v0_3 [3]), .B(
        MCInst1_MC3_v1_3 [3]), .Z(MCInst1_MC3_r3Inst_XORInst_0_3_n4 ) );
  AND2 FSMMUX_MUXInst_0_U3  ( .A(1'b1), .B(rst), .Z(FSMMUX_MUXInst_0_n1 ) );
  ORN2 FSMMUX_MUXInst_0_U2  ( .A(rst), .B(FSMUpdate[0]), .Z(
        FSMMUX_MUXInst_0_n2 ) );
  ORN2 FSMMUX_MUXInst_0_U1  ( .A(FSMMUX_MUXInst_0_n1 ), .B(
        FSMMUX_MUXInst_0_n2 ), .Z(FSMSelected[0]) );
  AND2 FSMMUX_MUXInst_1_U3  ( .A(1'b0), .B(rst), .Z(FSMMUX_MUXInst_1_n1 ) );
  ORN2 FSMMUX_MUXInst_1_U2  ( .A(rst), .B(FSMUpdate[1]), .Z(
        FSMMUX_MUXInst_1_n2 ) );
  ORN2 FSMMUX_MUXInst_1_U1  ( .A(FSMMUX_MUXInst_1_n1 ), .B(
        FSMMUX_MUXInst_1_n2 ), .Z(FSMSelected[1]) );
  AND2 FSMMUX_MUXInst_2_U3  ( .A(1'b0), .B(rst), .Z(FSMMUX_MUXInst_2_n1 ) );
  ORN2 FSMMUX_MUXInst_2_U2  ( .A(rst), .B(FSMUpdate[2]), .Z(
        FSMMUX_MUXInst_2_n2 ) );
  ORN2 FSMMUX_MUXInst_2_U1  ( .A(FSMMUX_MUXInst_2_n1 ), .B(
        FSMMUX_MUXInst_2_n2 ), .Z(FSMSelected[2]) );
  AND2 FSMMUX_MUXInst_3_U3  ( .A(1'b0), .B(rst), .Z(FSMMUX_MUXInst_3_n1 ) );
  ORN2 FSMMUX_MUXInst_3_U2  ( .A(rst), .B(FSMUpdate[3]), .Z(
        FSMMUX_MUXInst_3_n2 ) );
  ORN2 FSMMUX_MUXInst_3_U1  ( .A(FSMMUX_MUXInst_3_n1 ), .B(
        FSMMUX_MUXInst_3_n2 ), .Z(FSMSelected[3]) );
  AND2 FSMMUX_MUXInst_4_U3  ( .A(1'b0), .B(rst), .Z(FSMMUX_MUXInst_4_n1 ) );
  ORN2 FSMMUX_MUXInst_4_U2  ( .A(rst), .B(FSMUpdate[4]), .Z(
        FSMMUX_MUXInst_4_n2 ) );
  ORN2 FSMMUX_MUXInst_4_U1  ( .A(FSMMUX_MUXInst_4_n1 ), .B(
        FSMMUX_MUXInst_4_n2 ), .Z(FSMSelected[4]) );
  AND2 FSMMUX_MUXInst_5_U3  ( .A(1'b0), .B(rst), .Z(FSMMUX_MUXInst_5_n1 ) );
  ORN2 FSMMUX_MUXInst_5_U2  ( .A(rst), .B(FSMUpdate[5]), .Z(
        FSMMUX_MUXInst_5_n2 ) );
  ORN2 FSMMUX_MUXInst_5_U1  ( .A(FSMMUX_MUXInst_5_n1 ), .B(
        FSMMUX_MUXInst_5_n2 ), .Z(FSMSelected[5]) );
  DFF FSMReg_s_current_state_reg[0]  ( .D(FSMSelected[0]), .CP(clk), .Q(
        FSMUpdate[1]) );
  DFF FSMReg_s_current_state_reg[1]  ( .D(FSMSelected[1]), .CP(clk), .Q(
        FSM[1]) );
  DFF FSMReg_s_current_state_reg[2]  ( .D(FSMSelected[2]), .CP(clk), .Q(
        FSMUpdate[3]) );
  DFF FSMReg_s_current_state_reg[3]  ( .D(FSMSelected[3]), .CP(clk), .Q(
        FSMUpdate[4]) );
  DFF FSMReg_s_current_state_reg[4]  ( .D(FSMSelected[4]), .CP(clk), .Q(
        FSM[4]) );
  DFF FSMReg_s_current_state_reg[5]  ( .D(FSMSelected[5]), .CP(clk), .Q(
        FSM[5]) );
  AND2 FSMUpdateInst_StateUpdateInst_0_U7  ( .A(FSM[4]), .B(FSM[5]), .Z(
        FSMUpdateInst_StateUpdateInst_0_n1 ) );
  AND2 FSMUpdateInst_StateUpdateInst_0_U6  ( .A(FSM[1]), .B(FSMUpdate[1]), 
        .Z(FSMUpdateInst_StateUpdateInst_0_n5 ) );
  OR2 FSMUpdateInst_StateUpdateInst_0_U5  ( .A(FSMUpdate[4]), .B(FSMUpdate[3]), .Z(FSMUpdateInst_StateUpdateInst_0_n6 ) );
  BIC2 FSMUpdateInst_StateUpdateInst_0_U4  ( .A(
        FSMUpdateInst_StateUpdateInst_0_n5 ), .B(
        FSMUpdateInst_StateUpdateInst_0_n6 ), .Z(
        FSMUpdateInst_StateUpdateInst_0_n4 ) );
  ORN2 FSMUpdateInst_StateUpdateInst_0_U3  ( .A(
        FSMUpdateInst_StateUpdateInst_0_n4 ), .B(FSM[5]), .Z(
        FSMUpdateInst_StateUpdateInst_0_n3 ) );
  ORN2 FSMUpdateInst_StateUpdateInst_0_U2  ( .A(FSM[4]), .B(
        FSMUpdateInst_StateUpdateInst_0_n3 ), .Z(
        FSMUpdateInst_StateUpdateInst_0_n2 ) );
  ORN2 FSMUpdateInst_StateUpdateInst_0_U1  ( .A(
        FSMUpdateInst_StateUpdateInst_0_n1 ), .B(
        FSMUpdateInst_StateUpdateInst_0_n2 ), .Z(FSMUpdate[0]) );
  OR2 FSMUpdateInst_StateUpdateInst_2_U5  ( .A(FSM[4]), .B(FSMUpdate[4]), .Z(
        FSMUpdateInst_StateUpdateInst_2_n4 ) );
  OR2 FSMUpdateInst_StateUpdateInst_2_U4  ( .A(FSMUpdate[3]), .B(
        FSMUpdateInst_StateUpdateInst_2_n4 ), .Z(
        FSMUpdateInst_StateUpdateInst_2_n2 ) );
  AND2 FSMUpdateInst_StateUpdateInst_2_U3  ( .A(FSM[5]), .B(FSMUpdate[1]), 
        .Z(FSMUpdateInst_StateUpdateInst_2_n3 ) );
  ORN2 FSMUpdateInst_StateUpdateInst_2_U2  ( .A(
        FSMUpdateInst_StateUpdateInst_2_n2 ), .B(
        FSMUpdateInst_StateUpdateInst_2_n3 ), .Z(
        FSMUpdateInst_StateUpdateInst_2_n1 ) );
  AND2 FSMUpdateInst_StateUpdateInst_2_U1  ( .A(FSM[1]), .B(
        FSMUpdateInst_StateUpdateInst_2_n1 ), .Z(FSMUpdate[2]) );
  OR2 FSMUpdateInst_StateUpdateInst_5_U5  ( .A(FSMUpdate[4]), .B(FSMUpdate[3]), .Z(FSMUpdateInst_StateUpdateInst_5_n4 ) );
  ORN2 FSMUpdateInst_StateUpdateInst_5_U4  ( .A(
        FSMUpdateInst_StateUpdateInst_5_n4 ), .B(FSMUpdate[1]), .Z(
        FSMUpdateInst_StateUpdateInst_5_n2 ) );
  AND2 FSMUpdateInst_StateUpdateInst_5_U3  ( .A(FSM[5]), .B(FSM[1]), .Z(
        FSMUpdateInst_StateUpdateInst_5_n3 ) );
  ORN2 FSMUpdateInst_StateUpdateInst_5_U2  ( .A(
        FSMUpdateInst_StateUpdateInst_5_n2 ), .B(
        FSMUpdateInst_StateUpdateInst_5_n3 ), .Z(
        FSMUpdateInst_StateUpdateInst_5_n1 ) );
  ORN2 FSMUpdateInst_StateUpdateInst_5_U1  ( .A(FSM[4]), .B(
        FSMUpdateInst_StateUpdateInst_5_n1 ), .Z(FSMUpdate[5]) );
  ORN2 FSMSignalsInst_AddKeyInst_U15  ( .A(FSM[4]), .B(FSMUpdate[4]), .Z(
        FSMSignalsInst_AddKeyInst_n13 ) );
  ORN2 FSMSignalsInst_AddKeyInst_U14  ( .A(FSM[5]), .B(FSM[4]), .Z(
        FSMSignalsInst_AddKeyInst_n14 ) );
  AND2 FSMSignalsInst_AddKeyInst_U13  ( .A(FSMSignalsInst_AddKeyInst_n13 ), 
        .B(FSMSignalsInst_AddKeyInst_n14 ), .Z(
        FSMSignalsInst_AddKeyInst_n12 ) );
  BIC2 FSMSignalsInst_AddKeyInst_U12  ( .A(FSMSignalsInst_AddKeyInst_n12 ), 
        .B(FSM[1]), .Z(FSMSignalsInst_AddKeyInst_n11 ) );
  AND2 FSMSignalsInst_AddKeyInst_U11  ( .A(FSMSignalsInst_AddKeyInst_n11 ), 
        .B(FSMUpdate[1]), .Z(FSMSignalsInst_AddKeyInst_n10 ) );
  BIC2 FSMSignalsInst_AddKeyInst_U10  ( .A(FSMSignalsInst_AddKeyInst_n10 ), 
        .B(FSMUpdate[3]), .Z(FSMSignalsInst_AddKeyInst_n1 ) );
  BIC2 FSMSignalsInst_AddKeyInst_U9  ( .A(FSMUpdate[1]), .B(FSM[5]), .Z(
        FSMSignalsInst_AddKeyInst_n9 ) );
  ORN2 FSMSignalsInst_AddKeyInst_U8  ( .A(FSMSignalsInst_AddKeyInst_n9 ), 
        .B(FSMUpdate[4]), .Z(FSMSignalsInst_AddKeyInst_n5 ) );
  BIC2 FSMSignalsInst_AddKeyInst_U7  ( .A(FSM[5]), .B(FSMUpdate[1]), .Z(
        FSMSignalsInst_AddKeyInst_n8 ) );
  ORN2 FSMSignalsInst_AddKeyInst_U6  ( .A(FSMSignalsInst_AddKeyInst_n8 ), 
        .B(FSM[1]), .Z(FSMSignalsInst_AddKeyInst_n7 ) );
  ORN2 FSMSignalsInst_AddKeyInst_U5  ( .A(FSMUpdate[4]), .B(
        FSMSignalsInst_AddKeyInst_n7 ), .Z(FSMSignalsInst_AddKeyInst_n6 ) );
  AND2 FSMSignalsInst_AddKeyInst_U4  ( .A(FSMSignalsInst_AddKeyInst_n5 ), 
        .B(FSMSignalsInst_AddKeyInst_n6 ), .Z(FSMSignalsInst_AddKeyInst_n4 )
         );
  AND2 FSMSignalsInst_AddKeyInst_U3  ( .A(FSM[4]), .B(
        FSMSignalsInst_AddKeyInst_n4 ), .Z(FSMSignalsInst_AddKeyInst_n3 ) );
  AND2 FSMSignalsInst_AddKeyInst_U2  ( .A(FSMUpdate[3]), .B(
        FSMSignalsInst_AddKeyInst_n3 ), .Z(FSMSignalsInst_AddKeyInst_n2 ) );
  OR2 FSMSignalsInst_AddKeyInst_U1  ( .A(FSMSignalsInst_AddKeyInst_n1 ), .B(
        FSMSignalsInst_AddKeyInst_n2 ), .Z(AddKey) );
  AND2 FSMSignalsInst_doneInst_U5  ( .A(FSM[4]), .B(FSMUpdate[1]), .Z(
        FSMSignalsInst_doneInst_n4 ) );
  AND2 FSMSignalsInst_doneInst_U4  ( .A(FSMSignalsInst_doneInst_n4 ), .B(
        FSM[5]), .Z(FSMSignalsInst_doneInst_n1 ) );
  OR2 FSMSignalsInst_doneInst_U3  ( .A(FSMUpdate[4]), .B(FSMUpdate[3]), .Z(
        FSMSignalsInst_doneInst_n3 ) );
  OR2 FSMSignalsInst_doneInst_U2  ( .A(FSM[1]), .B(
        FSMSignalsInst_doneInst_n3 ), .Z(FSMSignalsInst_doneInst_n2 ) );
  BIC2 FSMSignalsInst_doneInst_U1  ( .A(FSMSignalsInst_doneInst_n1 ), .B(
        FSMSignalsInst_doneInst_n2 ), .Z(done) );
endmodule

